��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
�쬨����&}G�Bo�=�׎Z��1�� ��aC&}N��c��a)QP�2v�l��k�G� oF��T%���Z�]��c�ϏL��著3����Z��	s Pިw�]p���@Khy��Ɋ2���[�2M���q�Q�J��J�K�\����n}���:q�ֽ���ڵ&� ��t;��'��hD��دػ`�y��F����0��T&9���5�ۡ�q����a�i��
�D�J\˘K,DH~b�}�|�9Y--_LF�+$�0�"sux��a��q;�	K[nJE��Ȱ
0��o�rMٴ���	_���m��b�	؛A �oɔ���-�aw̫��s#�k�bUj>�_v�T	l+3]����o�@|�-�R��ʙ[
Xs�9� �[v7��t'|�"z�LeN��*��������\`hA'���h�����'J'b�@Vt��e�R;&Y�C;*�OղlH̰6;�X,j&3���%�`�����	���c6�;���	��z;��W���-).�hVۯ%���S�K7 ����M�fƏǝ��:�����a�E�8؞��t�����H�>����)�����	5���FӨ�.�Il�����G;c�O��<�b�l���u �o��R�%�)�Z������]������R����'4�F�t ��֌��{Z������mi��\P��_��!�/�����Ì�$��k ��F�ua^(��S[ezu�C��������F �}<��������C�d��а;�%�.�
�
���	]l������3�o~���v1�63J�E��	|�t)�����G+رT?C�K| Ư���	����7y�<�22N���K����Lt�OV�bbߣ:xg����N8���JRql�c"�|~��*��<k��w �	Z�Keq��ͥn���۩q�s��V5��r�Y�ZF_-
�.Q���&��g-_z�q��:�����b�a]�5�����C�4K�p��"���w��v�1��I�j�6�[�7[��LͬO"~�霍@�y�����I�"j�pz�Π�q�����H]ݥC�w�b�~&�hܟ-���Vbh��ܸ��+��=S�&���W� ����˩�[Q�yV32m$}�Rϩ�c�Cx4�VUs)�mT��zi��?��v�G[���\&�,h��\���䲣	U�BC�^;u�D|����^��*{��\�#��Nͣ���Z��X��݉��#�~���-Of|��{��;~�� �i��vf�4t�B�#�S�LT���w��'�΃��E&uWP�>���i�,X��t��4vD���Qo�Q��i):�߫�餝�k�c룯Ĕj�2��сS��X*�T��j�d�dF�5�՝��Z1��`F��.���,�U	Uk��Ų����D����yJ�N�'"��3�X�ն����dGx|tO��S���H��HpRe��(#Z��
��K�V���%jW�*6h`��QKRa����?���qb��̈w^����>/�gk2� �=!�\�ͱ��[r�6�Id�v\�A���B��4j�~Y#(h�bz;��֬��Yhh�}�'��ٙ-"? !n�>����t}�;?�m�l��M[�6��4R^ɞU��.0J5y���w	�����qÔP6R��,~0�:;�O�^2��ݐ����2�ѿ���Y���w��`�o���b���K�n{[�oK�O�����7�/$�wg}��R����[��[$p�8֗�Y�Z7�7�0��%��8�������d��F�#��T1���I�=;�l�3�k���S��e�4�����~;M�2����!"'RO0�-��B��?pЏ����[�ac��lO����&y��R�Cӯ��C4�[܂\��:�����G�Ƭb󁆠^��,7")��$Xp�mʋ�R,��cY6����4���#��K���ku����
��N�,��wI,)7L���A}��$��;<���EjY8ёw\���.�+�ω���������-�[lH�ρvE��