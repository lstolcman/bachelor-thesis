��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�O�5t�"��� ĸN�V�)Xq���!oA�㝣�V!��(r����6��DԓB�ee[�4���j#r٧a��������9��նwo6���6�"��ݿw�{,c�x���	��
`wgc���2�`t���o�(6Q�����w<�t��B�8�Q����/�=xy��@}W�U���9+�Х�4��@�L)���+�K��O�1��ºϷŷ�B&8�R6��Ե6t5�eD����+��)���!"�+E߷nld��\!������x��w�i<.s��mE��_��R'�[E`=
�����.�8\�Q2~���Z���T$�/)�u�&<9�0��}���Jo�i۔��<j��,��-��)P�0�4�0J�e��i�V�#P韉��������ɩ�Uo�M�+c}�F���� ��a0ZI�GDrؿ��x���9k�XEE�W�A/<eU���
�	O��)J�=�i�phRC����Ŋ�P�����G��ij������]֔�N��'��^Z˫m��`��g����^+�Y��`�F2grRM�P�������Cw�ᗜ�q�j���a{��d���i�Q��i�*
{f ��9]���5x��AO�[P#��h��v�2.�/���v���xN�˫�WضW�ڷ������"�mo}�!�r`!�%���UP�_��d�L-u5��:�>�Mfů�Mxn�v�G�G5��cK��I��@5P@OmV�p`�a~ek��l�7B_��ƺ/(�WBYN�]���Vx�%��V�z��H��2O�F,���������+
��l�HN�/V������C�odIB�~�2 �*d-w��N��T�8�I�욫��p��d�pߵgBq]H��@w���=�g�0���" <=���&I�恍5w�Z�M��.n�e=�i2�nL�H�!���eQGZtuRL�C�+�j��"%���N�	ۢBe^M�M^`��mb�]%�+��)	�Vb=9��a ���Dki�OV�P\O�n,-��C�z;9E_kOP���ޅP��J�n�.30���2���E�\���
��B��	J>b�
`��ő� V���V��$#�gOq@.�7�8|AtŜX����@�Wr����x��Tr٭��eW��vsO��С���(r%'�Ֆ����g�D�lw@ ��Y�p�&M^���O�#��D)	e��o��Y;ǌ�MFz�z�ē���.׼�t(�#j�9�����P8,�O�ѷ��i�q�$�.�LJv���s;��@�r�8\�0x�k��t@s���F8K�d�ܮ�/݊e�GEr%��(��'���z��ױ'��Ȧ���k-$��y���lr��a���8��/�N(+pZL<�M�z��k��[y�_��N�.���c{.���Q�U	a����&(�	)5��+\�;�u����`�������������])�t����n�b�%��ƅ��9�H�����1��΄є�ɾ�:��3"�9
�}\����&�@b� �~����#��w��Պ+C���h��'�	L;D�4��-��]�Г��D�2a��H��o�G���.X/�`�JH<�iWRvDE�]���"�Y�]������_ٌn�	|���݈���u]����4}�8�ɤ��h%!k�;���(�9�~�����w.4��`ش�;g�d?�iGx��o_�{^v=�ʪO:yi��e��5L�+f�څI �D����H-�8�ś6,t�� v�n3�g#�#a�#W�-��hU�-+������贝�n�5�*��eZ�R�ȋ�p^�G�n��:����{����g�ݵ��!�
0�U/���M�U=��?'��ZL��ŋ̗=�	�?U�f��)Ml���؊�r�ɚ!�4��5�����oB�'Hk6Uk��s��-�UE�YsD���N�\{�1_S�}_)�.�������ɂ�c��*��)�y��|'�k��S*��+i<��}/p<�|b���j�v ��2��z�%Tƹ��19U|Z~��7`Q���p�|�6��E�)�q`�Pe*J_���R �jk+t��Se�G��&��yK�i!r���o�&K/���][��5,�+��=ǎ�����7� ~��ž~��P�O冽A�
	�`S��R{"���o�pE#��_V�)M��,s��Dmĸ��E�`�[��#�W��/]r��ʏr�(X���ɅՄ��
.�֭�����Upz��ʥ��]t�����;��!7	�I�pǱ;v��e����m��Z�W�.!?r�� ��V�/g+��_[�݉����	�Z���*%��ŭN�Z�K��Y�>����RZ���G_2wg���#q
q�V۰��[E���.�Ϛv�K��������H�a�s}�%`�O=��snS���Ɲ���C��Ɋ�F�)ϝ=L��~��Y�q�d����wu}NߒHI��6�݈;RZ�'?�p8�I�@)������|�Xv	�q��+����s�a�����!�ji0�_�Y�JI\�����ݷ,�������
g+��<�^��S� ���Y�� k�A�7�����4=��+���pno�H^Ϳ��M��<�y#�ʝ;@q'�$r����k�X��`��	�$��^��~
(�H�9mݘ�7Z��0��ݞ��B�[�$\=�/� ��߮ē�;BH������&>IkL�l���  I!ɋa�'v��h��Tv¹Rew�����n�6λ0��z�Q= �p\oU�=
�E4�GP���h��s�wZ��jO-�=>�W���J���A�8b��wd�3T��G�Ymo�/��W�h�Ǌ$�vkA%/��	.�o��i>��p'Uݺl�1AL�B`���8�_گ�0�9�*ry1,ZQ�s�����ԫ-�Cb�`X������8J���uҽ��t6���hq�/�7��MPו���s�I*10/p$G��K��U*�f�R���K�?J�kj�Ũ���M)Lj��5����lV�`��a���� �{h;%�?kN�υئ�^p��p
��l��:a�fF��*\�����č»�+���G�3W���@�1g-\���I�ae~\렼��e{�����+��j�a�a�W�CV�Ơ��/������i��Ǘ���Iu{�R[�7z�(�q�c�V(7�y^�傩,n�X�x�%�( )����jj�?��j�A܎�n�/խ��aR
7�r��Ge���!�8�k��[������S9�V�IK~x�ql:�։��
�z%�l%�Ʉ+II�G r���R�3�A
�n�E�Il�wk�de\�3T�r����?Q>�iZ�1�B甆��(��٪Ux	Oj�$�Ğ����H!�vɦs)R*�~O��=|� B��z���A����\zUN��W4��&��|�`h���X�v�'1\@�<:w��.P_ 4jg\�sTQ�V�T�U������!73��4���6�F�y�aZ��_�7N����s�r�O�jR��f��D�b�2�Z����8	� r��SN�k�
[-�PX�e�~�8�U5�Z`Q=y������]?��A�t~==؂-�:���\Fg}�b���]]�BT�\�� #�ю2[����<O��׾�=�#$\V~�V��Xnjr~tTy�,���uc9��Cr������]�U�\���~l���F���n}�tՂ\�&�?� Эj�UU8�@�!��T�1���3�sA�
��з����V+�z`9eJ#���$� 
�6N��M/��D1,XzM�Dχ;�3�v�Õ���DA�hVH�<1��=ߊ�=��t�
�4d�=��3۰U�,����.���,t�.�m[�:\�4f��:��@���$7�xEFq������]���Ya��.(��f`����qm��ia��j�z���YL.��w�c���pY�N^�Y��Τ���H��kI���0�����䗗s>��h	�[{���y�5^:���NJ�f��*��,#�k����� (-\�RO*M3}Y� "��c�d��i��0G����#���������W��8aB>W_��-Y��l�Vs$ ɤJ�i8���g�Ӝ(�0P�v(��ö��UCNt�IP�d9Cڐ�� -�N����Z�d��C�s�T�lUq��(��&$�������
��)(`%2�96� 	�)�*8����n�ۍA���P���"��/�c�N-���+��Jϑ��h)e��n]zN+�",od�xU�0�#{�7�K�H�N!CA]�2�o.!��ws����q�k�_�t���I$K�\�����ȏ�t��V_�zY��	��:�҂�|�E��/Y���Hz,(0]S���lE��g1ؐ��Ro� ���hU�������yщ��v�li�3���O����'�c�¼��H�Rՠ�哛Kf� |I�מ�q�e%�
���"�m���}$_��j�>�]�T"�Ȃ�i;��	q*��ic_d�{D�9�T��-�z���b��^�ҭF|���:܀�0'(^��)(?���n�4r@�(b��*���y�ցW[�k���+͛`��8&#�Ӎ#���I`�� ZJZ�i�u�-߂?���N��_d�G�f8�IŎ��a�[�۩�j.��<��F�S	/�po:���`&<�\�p��X�{_*o���*�Iv��2<���,�#���?>�%�>������i���Y� ���Y�	N�]���HPi9����۠�0��¤��n��QK �[���C49��.wo�Ѝ���J>,����GO84��O�*XV��?�(�꾐��s�Hh�A�g�l�3�*tA��;E)��k����+��2��?w�t�]#ϕIpy�N����&A��*]�;0�������kĊ�E��RS-�.,�fܳv�s�m�G�-�U��<�����־�rh���z�x㳜�y���q�h�(Af�Ь~Sb�9�g��a�s84�uV/������0Su�@tE�����+�N�&ium��h�Ȓp������w�C�
"ф����P,�շr!D��%H>=�y߯z8� 7.c^���-g;�Лg��!�jV��� �s�b�0|����0�|�:�g��bڭk��yKl��7���m���Z2�i?��(0��;��ܗlI�)�.���N8	p���KT�9��
o��T(w�����ozl`DW_ϐp�*��jR�T�[$܇.�⋊�^�ɣ��?�yH+��#����n� (�Ox�-�2�����V��Q�N�u��^�oH(pć�P��N,)Y8�/�(F��n�O�%|�j��qڻH l�v��	L��K�X?�Z΢�����Y ;��_{�ޔ^����e��q����ѷ3�r��t�<RIm~֑��V#��x��̓��P�J�t�c�s,R���jz� ��;�	u�(�`X�6Ox�֒l��G1�eb$�������H��=���I�X 0<���x�O���K����L�v^(|��3�v;0l�'�ⶩ?	�+t��sqȩ�}8��{��`������ݻh�K���480f�?���(Z�Q]�l]����*��r�O��(3ғ)�r0� �۽ȑ�E�*'.n�����eaFr�A�Z��,,�M���p#�>X�
):��xaS�R!D��f����Hb�����'Û��	�@=0�<��rk�H�+����mG�J��1���(��0ȯ	/��>K/�ᔰg<�q�Xkj�V�ZŽ}J`!S���V��i'��=�	�ٴ-��#�lnl��t�<�mr�W����v믕�ϛ`DhQj��9yh¼�!0t/e%�OAq�;�䴱q�j5*��C�E���廁�5��?:����D�^�F����_'�ͥ1l��x4�����ɑ�*�cn��ً�;��VC�V��ب#��B�(��/9�/ok,H"7W?�������Y�$3����!�v�E�G q��M��*�qk<�	���w�{�����K$I͉4!���Oz�wh��iדD$A�~��۳ׅ~�S"+5��.�$!�˿sBb�R��n��L��t8�Cxfb#*��ԛp���WG��)����~e����D��*���[ǣ�^
�K=�>j��<��Cv�ƍ�S6��y�|8-���7h~Û]�������CPv�b!�~̲c�'�%/��X��<+&x���j�y��o�j�й^E9JLH���vЦشÜ�_mȮR%�D���O=�ʙvVؓpA~fV�َ��X�L���G�ny�}�b�zw~�T-)6�%F9��LZV�p��a���4��?x2T+b{�j�V����^m���xg�[�"�s}�p������A�3ͣ�<kڨC�Q�P]�
��c�Ð��uNOI3vGF���5���Os��~�ŔL9q����n����w��<�/r���AXj�
�i�Y�o�3�Z:�T�����m \Ҫ��m�ɛ��kOccS����i���A�����6N��(:�C0���qL2��c���,{M�L�W��*���8
���j��@.����Ct��]�������c�C��2�O��Ic��֙="��Q.t�[ƌ�/���N��or�ʰ���IVbx����P�8��w��9 �D�ߡ׹.*yc�4���E���x�h��΅���e���}|Z�|2a�(��q6��^#��M�ǰ�$�D����H��VC&y�q�M�a�8,c2n�G� [e�$<���b��E���}��N�gKT�������ⓟ��v�����֟|̞��Q��Ga�\���s��w����5�^��k;ʔ@�NHp���-��T( q��²�����Ӥ{D$��2�Zy�2iĔGg�&5��{Ď%�k� �k57������NKcf�]ĳ���U`��%'>�oNȔ��.S"���o��j�m'���F�� ^�+G�Y%���
����PJ��������0��'�_kP���}v��+Z#v�t���C�4w+N��ze���bj=�o�O	�%�n���}x�Jj8��[wߝ���-e;���$�}cX�����e��5���~�M7�n������wQ\�=`��_�4�bHqv��Cb�EkM`�N�E����K罠�;Q�N	�˘sB달,��>����˷���R�A��݊������U80[h�Al4>���ѫٱQV+��o��`��ܝ�)9���&1�(��Z�K.�p9�F��PF�!���
���Qo�퉎��Q�N-ӊ�C��9�aB`B4	��!/!:�l��5�3KPb9�w�q��L���n�O��;�#ȷV��3n2��������o�FEJb�s|R�cuI�x��?�5e��T8.�ݎ���8�%�F��1��`&J��h�z@�G��p+ʾ$kԨ^��C�@=n�P'�����Eƽ�تʿ��8� 8�s
�z�֔�Ç���v����ٟ�UY��ur$eu��t�f�;#>�3�v���}!�z�@��\(���V�nn۶s���;,W�s������/z�f�<�x�}T��ʉp���X��:C~PF3��.{��l)��3wO� T�/]�`*Ȅۅ̥���l��F1F��T��ui�$�,��qΖ��hs[�a�Rm��E�ː<���n�w�A�?���{`�F�v� ��mLQmgO��
ݱ����R�sdhGn�|�i�9a�\�>Rb*"2!ax�	׏�	ӱX[_#��JѦZ��=�QB�Si��+(ܕ$�`��"�W+_��(R�<^��,":�Ȱ�cUx;"�Q���!vE��+R�voj�t��ɟ�AR�����o����OF�w{c=7�1"�n�At
9�F��hT�]e:<x���^idH/8�w���w��tԓ�d��r�K��ҋ��	�MN�SE޿^���֍�����f�l�Z<�vb*HҌ>�Zhv��i�G�ND�]�-v*��G�h��9���b�����uM�E�oh�cq-��bBKa��5WF�Ys��K־}ﵥ�|wɖ����O� b�Jmc`���x6����%�ݞ�ڽQݠ4]�Faw$	��z�P���ٙ�NN�j3�b,�|I��wsW�n��ħ���v�F"鬯 ��^���U�ד�)o���͑5o�8��*v�T�U{"�A���IKf���=��:��?Lc�T��s)���-����*�s�5�?A_�E��ృ�c�g�����/z:'�����ƝQe����W������J�������gͩ��X�X����Jg��#����3킸�fЉ���L~v|<,�A`�L��:��Q' T�&��;��6!�^�޾�	/k���/�P�����L�2� h����#\��;	b������.�Q>�㕬�S��j��S#Tƥ�H@MN�'�FY�h�u��<��x'ޤ~Փ?�y�zX�p�^
��_�N��h�K�s�i.�.Nr1#��jJ﹩S�Z�͠"�U�%�����-�^�����$�p�k��{��������j�w�J8I1��m[�XB~J#��m���;q��w_{���ד�r�1����O�GP�J����v��>>q��M�4)����w�_ތ�R℻Xhs;�R�$6��E�υ�w��*ABgJ�Z��W��B�; �e����p ��VJ�`��1��	f��`�����BSYfL�����0�#C�4~�EF��C� +pu8?2��=�B/��Qj�d�����&1���$?q�?�g�.�$�$���)�L�-��w-���ܮ��'�Wi�Q��1�����gg��]x�T��`x8����@;&�)pA@Ԝ%����XKݏ��f��(���'޾�-r���]8'j���0i=[
\%c�����u��H�8a��š�����cj�1��&��\tI�Id"���\
�"])�?�O��*���\�5����-ƦCd*S����/>K�rhS�h5'�6�� C�D�aƕg�S�8� �
D��5��ص�x���y�^�L+������F�������n��������`�/�#���h�w���3�&/��!-�f�<��$�F���e���7e�n�LiU�,~��T�g;f��]O�r�~D�������/F{K�
Q�|����L��it�<�E8���D�@`�.�.�-4�1�0��>JD�ᕊ$js�Dn:��p�;�U?8�8�ᐞ���v�1�<Gܳ��d�1�6� (��d��S�T` �Ô(�$�%/c�i	�]�?�0�'z(2��K"��������uT^�3G��JB'%吢b�H[����O��SU��r��%	\��fে�2�d�;a�b�Y���~0q7��{}��ޫ��ZU���Ɔ��C�I�$�����<֓'`�O���b�F:��3�<J�o��qU{����
rtAˣ�^"�C�|,=f���:Y�-�S�E�z���<�yq_�;d/�b���v(H����n�h��b&]�H>��-�Gq�*O�b������k�u��+�������O����+��W��F��w�ϻ�"�Z:B_�U$�nЋ�⾵�<�Z=���$�M/ex�Z4������i���ܖ'��9ݽi��mn=,O7B�tti���4�̿.Y����l@��%+��&.�*y��$�'��!z��<��㠰]bo��{�M������f����,�A�D�1R�=�啙L���L�iZϋ10���r���
�I�� U�c7z�u��*3=��n��G?v L�HĚ%��T�Q��%t�~�^sy!��N�!��#S�`�����P�&�lL�y("��+�	M('�Qh5�kx�j��(3Mz)eo�i؜D���6oI�&�Tk{̈́�xX/l��z\��B^9:$l��i��hIlP5�6Ý��y�����XH�
CY!�S�3�m�n������ �
��+�|�$�"��$(��2O����'�@�'^i�<�:�R���oA���
���	�&����w�1��'CeeV��g8�}�
]84��h��W=�������I��q�z
�#�"���8Si��� U_&_��(�{j�/�X?��{��D��O?�Ԯ��Xa"����b�`ҙ�%ٝ/q_�kgka���(u�Zr��꼌������ ~�7�Gd�������t	JH�C���`�2��a�k�s�0S�ge����/�Bڇ�&[�B�^d�=H��4�a5DB>�2z�Y�׳~�����WV��m�@�c���q���/x	6�u�"ki���/4�(�K`�	��X�o��ve�������сYU6u��C�0�j��"�������
����,���`̀�<_��0
�d6� 0y ����!p�Ƅ1��
�B{�OF��,^���*��<tY|VG�x�X��&OX�m�ݒ〉+�s���T��ᖴ(��4�Y�/1��C�:��������6j =\}q�K&�%K���,����f��\i�z���X_��#PR~�U���&=�o��>���W���PÖ�����%�b�s}�T��1��F�5�/���i����>����,�Z�~������R9�ڈQJ���<����5ф�*Um���� 8�"�0�+���\��&uZ�R�h���kL��r��p�-.�[�ꊍf�"�������'l.5=?�V6p����fQ��6��ꤍM]��A!� ����TJ�>��� �p?P��n��
:R�'�:��
N�ޖf�]�Ċҗ�]���x�}�?���Ɨ�d~��]� ��v�K\�L�oB΋��u���W���O�\/�C�O�������	���q�bR g{���jaN/����`��#�� N#S��!2|�r�	[Cc�������J�0I2��\���μ^`�A=�@�����|�,7@��͢� ˽�zG��p�(m�}\�@Gn��w2��~��R����?bZ������a^s�H�y�K�h�$<����uv
��*H�~�[^-��͍��;������D�$���Ja�d� �ajO	�,�lmԯ'���g>q�{z,vJ�Qj6�����K1�;�Ca�Cw�70]**�R�	��C��{,e�gfr���]�c;m�x���*J�>m�@��l�:%	���MW�����<4饠qm�	̰O�0ppo���&�Cl�/� ӦK�� %��M����qk&��f� �� �}X=�_�$�zՙ��s�g�/�o�)���(�l����u�*τ����t��Iv��5C%��t�w4O�@�n�E<�3(u����Xy�O�MP�1�?�I⏳��nm�iQkU������Σ���y��p�&���y����e�TW�A��M�D"0r�ē����/[u��b�y�,�fH�.w���dr�[z5� �0��O��`~/��Z�"��U�9r��؂�k�t.�����BKr؊�����Q��+���z	�`���%�~�M� ��tߢ��߻L��~(��_�@ᙙ<�-�C'�)I��+W����Y����w�9�M���X���C"Y)Z;��v���>"~{T���Hѓ�������������Z����g|��w'���F��������x�/�����L9��U�9����i��^�;īA�_=T�W�4��([Z7tIA����Ҍ=�I6[+��6�ne��$9oQ ���8���;�=��W�`T�����,�릧*��nb�_YO&��ëz�&b��`�U�G�'�dyֿ��G�N�Z��"z����'��H<�� �w`�_u(\��6�q�|K�\��ZEn	�hE��A���i�?3 X�Ў�0�󏹭�X�ܢ�Yy�N�����hI򵘎��Y��GA��|��GR���1�c@��h2���Q� ���0ԇCB����P)�ۨ�<��l�f���й!Yo�uabx��DM�R�����(7UT~��l?��c������^�;����`ߤ� ��-!tu����
�����WQ��g����>��2Bl��26��}Vl�)z˾���r���(��/|�?�I|��L���2閉MZ�z���8O�ȑ�^b���ɦUK���.�AsG�r2-�c���C+"��z�p�&[7Ŏ�e@@PD����Lug핻��?vY=24�W�6V��dy�g���q��Ni����BY�I��/xԉ��!Il����"�����.qWE�S����д"65._�Z��4����G�I�}����.����~PԒ��%�A8����z�u�8��&#������$�zЧom�a�e��Vy_9����c'g�ܵ;0�T��4�év�� .f�g��%u5 5Es���4����t�����~�l��9�dMp��W~{V����_R�M��+$�-�h	����I�L�n�Im^��6�>o���b=�	ٞ0�b�t���A�N�:�=e���u������50
ra��C�ɓI�U��p �b�u��"����e�Qѳ�����ǅ�K2B� XH���e��aa-|�r��!��	��m���=�rМM����8�bo�rV�N�jMw�k��<�����W{����m:��{�!�`