��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6� '�7mF�Y��ߎ�~�+|���<�0g�s��\��[�� ~ ��a�j�}�T�X��: h��{o2]+�q?���Lo�c=i�$�^?���t�0I|4��(���������G�=�e��V��z�m��ٿ'�!Zd��������]?t��(�>ȣ�K�=�>>%`�8����8��kethq�����pb2E�fsV$ Ѱ��9����>�
Ls��W+�����0��$_�n��ܗ�՗��d;�Q�د�K��f����lm0}��	m��,y�����(�����\	�ї�S@5 �X/�ٞ����ǀH����*�o���D������
p���E����6��v�//���p(�w��wׄ.�6^�)��xy�p����g}9��l���ί��Mgò������ʝ��B���@���U�Exq�̼I%�%H_�J�DI�g�M����+NV��LK`����]�T�Ƒ�cu@�Ǭ�,�7 x�E�N�&�Pb��7���
��jL�&����\�S�<�e"R@ ��]���������Ȓ��:OT������oN+�;B�b
̸�E���@��D1�q���%��,m��gu?�g6�g�øZ���0�0�oRh:��Mk��YU77�bKj޼CV�a�ޅ{�H+*N��ts���l��d�j:_�V�`x=X��Z���F8���cɉ[&":����&4�dQ]�DI��g;W����������^�.�4ξ�'A�<�����A1�Y�\A���`�q�CQXk$>{�h��Ԧ,c�.	U.����] ���(�H/��+-����Z��jӏ9���9�t�̵'�8��q�[�Ұ6�c��a֜n��%��y/<�8ntʄ!����?ې�eq��QA�M���9�z�Č3�E8�������j��H&�M�W2�b�P��%r��b��s^�R�qHg�p����in�
�#�QqҞ"4����,��ʦ����,���t�\M�\I�����.X羃κ5`��~�  e8�)s=�{ܷ��|���mv7eG��z������:��qI�q�`�G�-T9�*r��Y9 oW�5x]�>�7i�*%�X��������