��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#��^��B�J��J�+.�&
\���S�%�eV�7������0g�{��c��0�Bз�;����{�_]<ym�nU"��5K�4j��ǽ�������X�n;��ݣ3A�ځY���}hXu*����8T��-��Ĝ׸��1�L�Fp5���8\���;��^D�����j�16�B>ƀو`���
@wrQ@�X���\��`z�k&ޥ����F�>�n/r���yE=��	�M�´Y�V��t�ME���T�VY��)ڪC�/��i�>�k)G(��T,�����	�,P�%�0|(��<���D�0��#�+�ᓇ�w!�v���g)Oi�-�o��͆�cCÎ�� �Ｗxܼ����AD�e�1��Q��嗨���<[W�k�5��>��#��N��>s�6N�g�����;rGXÃQH؀�o�CY���?����ݳ��G��b���y��i��<;��0T�}neGM�,�R���A��)/=�D*p��2��|D�m+^���M���1� Zvԇ[%�Q|fVN���x������WZ��C	Ip&��cD�߀�S�o>2T�e��-&���Iv����E�h2���:�n� �Zl��<��~%��dX��AL�r��{��u��,V{@+Q�:�@xQѯX�E���0;�Lwɵ��8xd����d��+�@ E1�3j�`HE<jX��?�\e�h���S�I�����[?jE������}B�:6u%�j�ߒ�9j��'y+�B�F�n.G���ۑU��|/�!�CP)S���֐�)q\o�{V��H0 i9���mC�kj�g.��]��(���2�O��5eHV��/�ݩo*���$�4��:��xf�F���
�n�����
��/a�{��������Zt�8�3��ز����L��0��pײ��,��9
�>ۉ�B��sx����n��DTA��{0��s�Do��}���>V��j���a���(���§Ҩ�|҂�z#�v����� ݇&���P��UsM�$��G���C+�ޚ�-�Kzh2b�\�[������TU��I��nau�"ho*�_^���?Ȭ.�K.�Q��5c�F��C6��bF����jU�6z�����A|�{흹Ǖ�W&�tޒ��!��>7��}#c����$#'n���7���L8�����O�kS�8�2��3f+Xx{u=��\��Qs�a�A�n��&��iU�a��U>u��֝��}��H��rv\IR�f�I8.��7r�N���z�_QP�4/�.(e�O����X1��fV/�f/_�D|FSL�]`�/�p�Jc&��[���JI�Zg�	�0�,��T*R�8ZT&�(�š�y���ž:���-��t�lˍ�3��D�����Sb
E�n5U2����
B0[r��w1��Vsb)��J���.�������������Y�ؔ~V������80�^$A��m^�E�;��b}��4\fh�(�����E�HÏ�a����� ٷAw��F��(k+��:�灴�9�^�i��