// megafunction wizard: %FIR II v15.1%
// GENERATION: XML
// fir_first.v

// Generated using ACDS version 15.1 185

`timescale 1 ps / 1 ps
module fir_first (
		input  wire        clk,              //                     clk.clk
		input  wire        reset_n,          //                     rst.reset_n
		input  wire [15:0] ast_sink_data,    //   avalon_streaming_sink.data
		input  wire        ast_sink_valid,   //                        .valid
		input  wire [1:0]  ast_sink_error,   //                        .error
		output wire [25:0] ast_source_data,  // avalon_streaming_source.data
		output wire        ast_source_valid, //                        .valid
		output wire [1:0]  ast_source_error  //                        .error
	);

	fir_first_0002 fir_first_inst (
		.clk              (clk),              //                     clk.clk
		.reset_n          (reset_n),          //                     rst.reset_n
		.ast_sink_data    (ast_sink_data),    //   avalon_streaming_sink.data
		.ast_sink_valid   (ast_sink_valid),   //                        .valid
		.ast_sink_error   (ast_sink_error),   //                        .error
		.ast_source_data  (ast_source_data),  // avalon_streaming_source.data
		.ast_source_valid (ast_source_valid), //                        .valid
		.ast_source_error (ast_source_error)  //                        .error
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2016 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_fir_compiler_ii" version="15.1" >
// Retrieval info: 	<generic name="filterType" value="decim" />
// Retrieval info: 	<generic name="interpFactor" value="1" />
// Retrieval info: 	<generic name="decimFactor" value="100" />
// Retrieval info: 	<generic name="symmetryMode" value="sym" />
// Retrieval info: 	<generic name="L_bandsFilter" value="1" />
// Retrieval info: 	<generic name="inputChannelNum" value="1" />
// Retrieval info: 	<generic name="clockRate" value="130" />
// Retrieval info: 	<generic name="clockSlack" value="0" />
// Retrieval info: 	<generic name="inputRate" value="130" />
// Retrieval info: 	<generic name="coeffReload" value="false" />
// Retrieval info: 	<generic name="baseAddress" value="0" />
// Retrieval info: 	<generic name="readWriteMode" value="read_write" />
// Retrieval info: 	<generic name="backPressure" value="false" />
// Retrieval info: 	<generic name="deviceFamily" value="Cyclone IV E" />
// Retrieval info: 	<generic name="speedGrade" value="fast" />
// Retrieval info: 	<generic name="delayRAMBlockThreshold" value="20" />
// Retrieval info: 	<generic name="dualMemDistRAMThreshold" value="1280" />
// Retrieval info: 	<generic name="mRAMThreshold" value="1000000" />
// Retrieval info: 	<generic name="hardMultiplierThreshold" value="-1" />
// Retrieval info: 	<generic name="reconfigurable" value="false" />
// Retrieval info: 	<generic name="num_modes" value="2" />
// Retrieval info: 	<generic name="reconfigurable_list" value="0" />
// Retrieval info: 	<generic name="MODE_STRING" value="None Set" />
// Retrieval info: 	<generic name="channelModes" value="0,1,2,3" />
// Retrieval info: 	<generic name="inputType" value="int" />
// Retrieval info: 	<generic name="inputBitWidth" value="16" />
// Retrieval info: 	<generic name="inputFracBitWidth" value="0" />
// Retrieval info: 	<generic name="coeffSetRealValue" value="1.57159478763E-7,9.91121276743E-8,3.46590455053E-8,-3.62938071403E-8,-1.13815267335E-7,-1.97947582979E-7,-2.8870508264E-7,-3.86072909296E-7,-4.90005825131E-7,-6.0042709453E-7,-7.17227452294E-7,-8.40264164012E-7,-9.69360185384E-7,-1.10430342711E-6,-1.24484613176E-6,-1.39070436888E-6,-1.54155765411E-6,-1.69704869824E-6,-1.85678329124E-6,-2.02033032645E-6,-2.18722196949E-6,-2.3569539761E-6,-2.5289861627E-6,-2.70274303305E-6,-2.87761456376E-6,-3.05295715119E-6,-3.22809472133E-6,-3.40232000421E-6,-3.57489597332E-6,-3.74505745035E-6,-3.91201287466E-6,-4.07494623652E-6,-4.23301917224E-6,-4.38537321903E-6,-4.53113222638E-6,-4.66940492044E-6,-4.79928761706E-6,-4.91986707837E-6,-5.03022350738E-6,-5.12943367417E-6,-5.21657416674E-6,-5.29072475882E-6,-5.35097188638E-6,-5.39641222386E-6,-5.42615635069E-6,-5.43933249769E-6,-5.43509036295E-6,-5.41260498556E-6,-5.37108066552E-6,-5.30975491746E-6,-5.22790244519E-6,-5.12483912398E-6,-4.99992597666E-6,-4.85257312951E-6,-4.68224373357E-6,-4.48845783642E-6,-4.27079618962E-6,-4.02890397645E-6,-3.76249444454E-6,-3.47135242796E-6,-3.15533774304E-6,-2.81438844241E-6,-2.44852391163E-6,-2.05784779281E-6,-1.64255072004E-6,-1.20291285131E-6,-7.39306182039E-7,-2.52196625692E-7,2.57854152898E-7,7.9018716518E-7,1.3440448009E-6,1.91856981725E-6,2.51280462732E-6,3.12569089944E-6,3.75606947807E-6,4.40268063655E-6,5.06416467064E-6,5.73906284141E-6,6.42581867484E-6,7.12277962456E-6,7.82819910319E-6,8.54023888662E-6,9.25697189459E-6,9.97638534947E-6,1.06963843144E-5,1.14147956104E-5,1.21293721108E-5,1.28377974104E-5,1.35376908648E-5,1.42266129954E-5,1.49020712518E-5,1.55615261255E-5,1.62023976024E-5,1.68220719474E-5,1.74179088046E-5,1.79872486024E-5,1.8527420248E-5,1.90357490935E-5,1.95095651587E-5,1.99462115893E-5,2.03430533315E-5,2.0697486002E-5,2.10069449294E-5,2.12689143453E-5,2.14809366981E-5,2.16406220655E-5,2.17456576376E-5,2.17938172433E-5,2.17829708912E-5,2.17110942957E-5,2.15762783572E-5,2.1376738567E-5,2.11108243043E-5,2.07770279935E-5,2.037399409E-5,1.99005278608E-5,1.9355603929E-5,1.87383745463E-5,1.80481775635E-5,1.72845440642E-5,1.64472056296E-5,1.55361012017E-5,1.4551383514E-5,1.34934250561E-5,1.23628235441E-5,1.11604068639E-5,9.88723746091E-6,8.54461614496E-6,7.13408528618E-6,5.65743137357E-6,4.11668691268E-6,2.51413163881E-6,8.52293023823E-7,-8.66053943434E-7,-2.63788772171E-6,-4.45994194356E-6,-6.32870791796E-6,-8.24043792207E-6,-1.01911492929E-5,-1.21766293272E-5,-1.41924409966E-5,-1.62339294804E-5,-1.82962295197E-5,-2.03742735901E-5,-2.24628008913E-5,-2.45563671463E-5,-2.66493552025E-5,-2.87359864236E-5,-3.0810332859E-5,-3.28663301729E-5,-3.48977913156E-5,-3.68984209147E-5,-3.88618303614E-5,-4.07815535658E-5,-4.26510633501E-5,-4.44637884491E-5,-4.62131310815E-5,-4.78924850557E-5,-4.94952543694E-5,-5.10148722617E-5,-5.24448206717E-5,-5.37786500578E-5,-5.50099995284E-5,-5.61326172323E-5,-5.71403809565E-5,-5.80273188753E-5,-5.87876303958E-5,-5.94157070391E-5,-5.99061533E-5,-6.02538074218E-5,-6.04537620253E-5,-6.05013845288E-5,-6.03923372942E-5,-6.01225974348E-5,-5.96884762194E-5,-5.90866380079E-5,-5.83141186509E-5,-5.73683432897E-5,-5.62471434896E-5,-5.49487736423E-5,-5.34719265734E-5,-5.18157482904E-5,-4.99798518098E-5,-4.7964330002E-5,-4.57697673941E-5,-4.33972508717E-5,-4.08483792261E-5,-3.81252714894E-5,-3.52305740093E-5,-3.21674662109E-5,-2.89396650019E-5,-2.55514277751E-5,-2.20075539692E-5,-1.83133851494E-5,-1.4474803574E-5,-1.04982292173E-5,-6.39061522084E-6,-2.1594417515E-6,2.18729175344E-6,6.64107596782E-6,1.11929026956E-5,1.58332775328E-5,2.05522341735E-5,2.53393503567E-5,3.01837654462E-5,3.50741996291E-5,3.99989747174E-5,4.49460365274E-5,4.99029788116E-5,5.4857068708E-5,5.97952736713E-5,6.47042898419E-5,6.95705718058E-5,7.43803636921E-5,7.91197315517E-5,8.37745969544E-5,8.83307717371E-5,9.27739938321E-5,9.7089964099E-5,1.0126438408E-4,1.05282994593E-4,1.09131615075E-4,1.12796183583E-4,1.1626279735E-4,1.19517753808E-4,1.22547591964E-4,1.25339134021E-4,1.2787952715E-4,1.30156285279E-4,1.32157330805E-4,1.33871036094E-4,1.35286264666E-4,1.36392411938E-4,1.37179445401E-4,1.37637944116E-4,1.37759137404E-4,1.37534942599E-4,1.36958001758E-4,1.36021717192E-4,1.34720285698E-4,1.33048731378E-4,1.31002936925E-4,1.28579673251E-4,1.25776627354E-4,1.22592428301E-4,1.19026671229E-4,1.15079939246E-4,1.10753823145E-4,1.06050938809E-4,1.0097494225E-4,9.55305421482E-5,8.97235098509E-5,8.35606867176E-5,7.70499887611E-5,7.0200408507E-5,6.3022014014E-5,5.55259450006E-5,4.77244060316E-5,3.96306567229E-5,3.12589989342E-5,2.26247609219E-5,1.3744278437E-5,4.63487275692E-6,-4.68517434806E-6,-1.41966487088E-5,-2.38794348944E-5,-3.37125503693E-5,-4.36741826375E-5,-5.37417293322E-5,-6.38918412007E-5,-7.41004679264E-5,-8.43429067189E-5,-9.45938535969E-5,-1.04827457278E-4,-1.1501737558E-4,-1.2513683424E-4,-1.35158688023E-4,-1.45055484021E-4,-1.54799527004E-4,-1.64362946688E-4,-1.73717766784E-4,-1.8283597567E-4,-1.91689598536E-4,-2.00250770834E-4,-2.08491812867E-4,-2.1638530533E-4,-2.23904165635E-4,-2.31021724825E-4,-2.37711804881E-4,-2.43948796229E-4,-2.49707735249E-4,-2.54964381576E-4,-2.59695294983E-4,-2.63877911642E-4,-2.67490619546E-4,-2.70512832876E-4,-2.72925065104E-4,-2.74709000611E-4,-2.75847564599E-4,-2.76324991098E-4,-2.76126888837E-4,-2.75240304773E-4,-2.73653785081E-4,-2.71357433368E-4,-2.68342965946E-4,-2.64603763935E-4,-2.60134922016E-4,-2.54933293648E-4,-2.48997532554E-4,-2.42328130319E-4,-2.3492744991E-4,-2.26799754982E-4,-2.17951234788E-4,-2.08390024582E-4,-1.98126221357E-4,-1.87171894801E-4,-1.75541093365E-4,-1.63249845326E-4,-1.50316154769E-4,-1.36759992395E-4,-1.22603281097E-4,-1.07869876246E-4,-9.2585540638E-5,-7.67779140932E-5,-6.04764776647E-5,-4.37125124789E-5,-2.65190532073E-5,-8.93083620082E-6,9.01575767296E-6,2.72827654338E-5,4.58307095641E-5,6.46186706703E-5,8.36043651309E-5,1.02744227618E-4,1.21993498359E-4,1.41306315006E-4,1.60635808941E-4,1.79934205856E-4,1.9915293042E-4,2.1824271483E-4,2.37153711042E-4,2.55835606441E-4,2.74237742731E-4,2.92309237782E-4,3.09999110175E-4,3.27256406169E-4,3.44030328815E-4,3.60270368914E-4,3.7592643751E-4,3.90948999631E-4,4.05289208918E-4,4.18899042855E-4,4.31731438225E-4,4.43740426488E-4,4.54881268705E-4,4.65110589675E-4,4.74386510919E-4,4.82668782164E-4,4.89918910958E-4,4.96100290064E-4,5.01178322269E-4,5.05120542245E-4,5.07896735112E-4,5.09479051343E-4,5.09842117659E-4,5.08963143575E-4,5.06822023246E-4,5.03401432282E-4,4.98686919215E-4,4.92666991278E-4,4.85333194213E-4,4.76680185787E-4,4.66705802747E-4,4.55411120919E-4,4.42800508207E-4,4.2888167024E-4,4.13665688416E-4,3.97167050157E-4,3.79403671136E-4,3.60396909327E-4,3.40171570685E-4,3.18755906318E-4,2.96181601028E-4,2.72483753092E-4,2.47700845219E-4,2.21874706598E-4,1.95050465988E-4,1.67276495838E-4,1.38604347426E-4,1.09088677034E-4,7.87871632007E-5,4.77604151312E-5,1.6071872327E-5,-1.62123044304E-5,-4.90233506197E-5,-8.22900238827E-5,-1.15938738109E-4,-1.49893705498E-4,-1.84077086373E-4,-2.18409146495E-4,-2.52808421608E-4,-2.87191888921E-4,-3.21475145202E-4,-3.55572591167E-4,-3.89397621785E-4,-4.2286282214E-4,-4.55880168442E-4,-4.88361233775E-4,-5.2021739815E-4,-5.51360062419E-4,-5.81700865572E-4,-6.11151904944E-4,-6.39625958839E-4,-6.67036711053E-4,-6.93298976788E-4,-7.18328929418E-4,-7.4204432756E-4,-7.64364741917E-4,-7.85211781324E-4,-8.04509317428E-4,-8.22183707452E-4,-8.38164014458E-4,-8.52382224533E-4,-8.64773460339E-4,-8.75276190437E-4,-8.83832433818E-4,-8.90387959083E-4,-8.94892477691E-4,-8.97299830737E-4,-8.97568168691E-4,-8.95660123576E-4,-8.91542973049E-4,-8.85188795861E-4,-8.76574618204E-4,-8.65682550454E-4,-8.52499913825E-4,-8.37019356503E-4,-8.19238958798E-4,-7.99162326919E-4,-7.76798674973E-4,-7.52162894803E-4,-7.25275613347E-4,-6.96163237162E-4,-6.64857983845E-4,-6.31397900065E-4,-5.95826865982E-4,-5.58194585818E-4,-5.18556564426E-4,-4.76974069687E-4,-4.33514080627E-4,-3.88249221164E-4,-3.41257679427E-4,-2.92623112641E-4,-2.42434537577E-4,-1.9078620662E-4,-1.37777469543E-4,-8.35126210986E-5,-2.81007345821E-5,2.83445184444E-5,8.57050620473E-5,1.43858623176E-4,2.02678951985E-4,2.62036054903E-4,3.21796440073E-4,3.81823374792E-4,4.41977154499E-4,5.02115382871E-4,5.62093262522E-4,6.21763895791E-4,6.80978595064E-4,7.39587202041E-4,7.97438415356E-4,8.54380125888E-4,9.10259759121E-4,9.64924623863E-4,0.00101822226659,0.00107000083074,0.0011201094201,0.00116839846563,0.00121472009489,0.00125892850323,0.00130088032593,0.00134043501055,0.0013774551885,0.00141180704517,0.00144336068749,0.0014719905084,0.00149757554702,0.00151999984396,0.00153915279069,0.00155492947218,0.00156723100198,0.0015759648489,0.00158104515433,0.00158239303956,0.00157993690213,0.00157361270043,0.0015633642259,0.00154914336189,0.00153091032849,0.00150863391272,0.00148229168325,0.00145187018899,0.00141736514104,0.0013787815772,0.00133613400864,0.0012894465481,0.00123875301903,0.00118409704541,0.00112553212163,0.00106312166208,9.96939030167E-4,9.27067546337E-4,8.53600474933E-4,7.76640989598E-4,6.96302117069E-4,6.12706659227E-4,5.25987093307E-4,4.36285450233E-4,3.43753171088E-4,2.4855094176E-4,1.50848505886E-4,5.08244562326E-5,-5.13339952819E-5,-1.55431268673E-4,-2.61263687788E-4,-3.68619772669E-4,-4.77280551986E-4,-5.87019895101E-4,-6.9760486327E-4,-8.08796079448E-4,-9.20348116129E-4,-0.00103200990057,-0.00114352513677,-0.00125463274344,-0.00136506730725,-0.00147455955058,-0.00158283681289,-0.00168962354485,-0.00179464181438,-0.0018976118236,-0.00199825243581,-0.00209628171133,-0.0021914174514,-0.00228337774888,-0.00237188154487,-0.00245664918993,-0.00253740300897,-0.00261386786864,-0.00268577174595,-0.00275284629712,-0.00281482742536,-0.00287145584653,-0.00292247765134,-0.00296764486305,-0.00300671598941,-0.00303945656762,-0.00306563970125,-0.00308504658786,-0.00309746703616,-0.00310269997161,-0.0031005539293,-0.00309084753302,-0.00307340995941,-0.0030480813861,-0.00301471342286,-0.00297316952474,-0.00292332538611,-0.00286506931481,-0.00279830258537,-0.0027229397705,-0.00263890904998,-0.0025461524961,-0.00244462633505,-0.00233430118339,-0.00221516225901,-0.00208720956602,-0.00195045805284,-0.00180493774325,-0.00165069383966,-0.0014877867984,-0.00131629237656,-0.00113630165023,-9.47921003712E-4,-7.5127208976E-4,-5.46491760512E-4,-3.33731969247E-4,-1.13159642847E-4,1.15043474904E-4,3.50681009077E-4,5.93542168231E-4,8.43401987657E-4,0.00110002160093,0.00136314853942,0.00163251705929,0.00190784849555,0.00218885164257,0.00247522316054,0.00276664800702,0.00306279989319,0.00336334176369,0.0036679262995,0.00397619644282,0.00428778594317,0.00460231992358,0.00491941546606,0.00523868221513,0.00555972299841,0.00588213446311,0.00620550772724,0.00652942904438,0.00685348048071,0.00717724060307,0.00750028517679,0.00782218787192,0.00814252097653,0.00846085611578,0.00877676497531,0.00908982002756,0.00939959525982,0.00970566690223,0.0100076141547,0.0103050199113,0.01059747148,0.010884561298,0.011165887639,0.0114410553133,0.0117096763576,0.0119713707141,0.0122257668972,0.0124725026467,0.0127112255661,0.0129415937445,0.0131632763615,0.0133759542729,0.0135793205774,0.0137730811617,0.0139569552241,0.014130675775,0.0142939901128,0.014446660276,0.0145884634682,0.0147191924573,0.0148386559466,0.0149466789178,0.0150431029453,0.0151277864804,0.0152006051059,0.0152614517597,0.0153102369275,0.0153468888035,0.01537135342,0.0153835947445,0.0153835947445,0.01537135342,0.0153468888035,0.0153102369275,0.0152614517597,0.0152006051059,0.0151277864804,0.0150431029453,0.0149466789178,0.0148386559466,0.0147191924573,0.0145884634682,0.014446660276,0.0142939901128,0.014130675775,0.0139569552241,0.0137730811617,0.0135793205774,0.0133759542729,0.0131632763615,0.0129415937445,0.0127112255661,0.0124725026467,0.0122257668972,0.0119713707141,0.0117096763576,0.0114410553133,0.011165887639,0.010884561298,0.01059747148,0.0103050199113,0.0100076141547,0.00970566690223,0.00939959525982,0.00908982002756,0.00877676497531,0.00846085611578,0.00814252097653,0.00782218787192,0.00750028517679,0.00717724060307,0.00685348048071,0.00652942904438,0.00620550772724,0.00588213446311,0.00555972299841,0.00523868221513,0.00491941546606,0.00460231992358,0.00428778594317,0.00397619644282,0.0036679262995,0.00336334176369,0.00306279989319,0.00276664800702,0.00247522316054,0.00218885164257,0.00190784849555,0.00163251705929,0.00136314853942,0.00110002160093,8.43401987657E-4,5.93542168231E-4,3.50681009077E-4,1.15043474904E-4,-1.13159642847E-4,-3.33731969247E-4,-5.46491760512E-4,-7.5127208976E-4,-9.47921003712E-4,-0.00113630165023,-0.00131629237656,-0.0014877867984,-0.00165069383966,-0.00180493774325,-0.00195045805284,-0.00208720956602,-0.00221516225901,-0.00233430118339,-0.00244462633505,-0.0025461524961,-0.00263890904998,-0.0027229397705,-0.00279830258537,-0.00286506931481,-0.00292332538611,-0.00297316952474,-0.00301471342286,-0.0030480813861,-0.00307340995941,-0.00309084753302,-0.0031005539293,-0.00310269997161,-0.00309746703616,-0.00308504658786,-0.00306563970125,-0.00303945656762,-0.00300671598941,-0.00296764486305,-0.00292247765134,-0.00287145584653,-0.00281482742536,-0.00275284629712,-0.00268577174595,-0.00261386786864,-0.00253740300897,-0.00245664918993,-0.00237188154487,-0.00228337774888,-0.0021914174514,-0.00209628171133,-0.00199825243581,-0.0018976118236,-0.00179464181438,-0.00168962354485,-0.00158283681289,-0.00147455955058,-0.00136506730725,-0.00125463274344,-0.00114352513677,-0.00103200990057,-9.20348116129E-4,-8.08796079448E-4,-6.9760486327E-4,-5.87019895101E-4,-4.77280551986E-4,-3.68619772669E-4,-2.61263687788E-4,-1.55431268673E-4,-5.13339952819E-5,5.08244562326E-5,1.50848505886E-4,2.4855094176E-4,3.43753171088E-4,4.36285450233E-4,5.25987093307E-4,6.12706659227E-4,6.96302117069E-4,7.76640989598E-4,8.53600474933E-4,9.27067546337E-4,9.96939030167E-4,0.00106312166208,0.00112553212163,0.00118409704541,0.00123875301903,0.0012894465481,0.00133613400864,0.0013787815772,0.00141736514104,0.00145187018899,0.00148229168325,0.00150863391272,0.00153091032849,0.00154914336189,0.0015633642259,0.00157361270043,0.00157993690213,0.00158239303956,0.00158104515433,0.0015759648489,0.00156723100198,0.00155492947218,0.00153915279069,0.00151999984396,0.00149757554702,0.0014719905084,0.00144336068749,0.00141180704517,0.0013774551885,0.00134043501055,0.00130088032593,0.00125892850323,0.00121472009489,0.00116839846563,0.0011201094201,0.00107000083074,0.00101822226659,9.64924623863E-4,9.10259759121E-4,8.54380125888E-4,7.97438415356E-4,7.39587202041E-4,6.80978595064E-4,6.21763895791E-4,5.62093262522E-4,5.02115382871E-4,4.41977154499E-4,3.81823374792E-4,3.21796440073E-4,2.62036054903E-4,2.02678951985E-4,1.43858623176E-4,8.57050620473E-5,2.83445184444E-5,-2.81007345821E-5,-8.35126210986E-5,-1.37777469543E-4,-1.9078620662E-4,-2.42434537577E-4,-2.92623112641E-4,-3.41257679427E-4,-3.88249221164E-4,-4.33514080627E-4,-4.76974069687E-4,-5.18556564426E-4,-5.58194585818E-4,-5.95826865982E-4,-6.31397900065E-4,-6.64857983845E-4,-6.96163237162E-4,-7.25275613347E-4,-7.52162894803E-4,-7.76798674973E-4,-7.99162326919E-4,-8.19238958798E-4,-8.37019356503E-4,-8.52499913825E-4,-8.65682550454E-4,-8.76574618204E-4,-8.85188795861E-4,-8.91542973049E-4,-8.95660123576E-4,-8.97568168691E-4,-8.97299830737E-4,-8.94892477691E-4,-8.90387959083E-4,-8.83832433818E-4,-8.75276190437E-4,-8.64773460339E-4,-8.52382224533E-4,-8.38164014458E-4,-8.22183707452E-4,-8.04509317428E-4,-7.85211781324E-4,-7.64364741917E-4,-7.4204432756E-4,-7.18328929418E-4,-6.93298976788E-4,-6.67036711053E-4,-6.39625958839E-4,-6.11151904944E-4,-5.81700865572E-4,-5.51360062419E-4,-5.2021739815E-4,-4.88361233775E-4,-4.55880168442E-4,-4.2286282214E-4,-3.89397621785E-4,-3.55572591167E-4,-3.21475145202E-4,-2.87191888921E-4,-2.52808421608E-4,-2.18409146495E-4,-1.84077086373E-4,-1.49893705498E-4,-1.15938738109E-4,-8.22900238827E-5,-4.90233506197E-5,-1.62123044304E-5,1.6071872327E-5,4.77604151312E-5,7.87871632007E-5,1.09088677034E-4,1.38604347426E-4,1.67276495838E-4,1.95050465988E-4,2.21874706598E-4,2.47700845219E-4,2.72483753092E-4,2.96181601028E-4,3.18755906318E-4,3.40171570685E-4,3.60396909327E-4,3.79403671136E-4,3.97167050157E-4,4.13665688416E-4,4.2888167024E-4,4.42800508207E-4,4.55411120919E-4,4.66705802747E-4,4.76680185787E-4,4.85333194213E-4,4.92666991278E-4,4.98686919215E-4,5.03401432282E-4,5.06822023246E-4,5.08963143575E-4,5.09842117659E-4,5.09479051343E-4,5.07896735112E-4,5.05120542245E-4,5.01178322269E-4,4.96100290064E-4,4.89918910958E-4,4.82668782164E-4,4.74386510919E-4,4.65110589675E-4,4.54881268705E-4,4.43740426488E-4,4.31731438225E-4,4.18899042855E-4,4.05289208918E-4,3.90948999631E-4,3.7592643751E-4,3.60270368914E-4,3.44030328815E-4,3.27256406169E-4,3.09999110175E-4,2.92309237782E-4,2.74237742731E-4,2.55835606441E-4,2.37153711042E-4,2.1824271483E-4,1.9915293042E-4,1.79934205856E-4,1.60635808941E-4,1.41306315006E-4,1.21993498359E-4,1.02744227618E-4,8.36043651309E-5,6.46186706703E-5,4.58307095641E-5,2.72827654338E-5,9.01575767296E-6,-8.93083620082E-6,-2.65190532073E-5,-4.37125124789E-5,-6.04764776647E-5,-7.67779140932E-5,-9.2585540638E-5,-1.07869876246E-4,-1.22603281097E-4,-1.36759992395E-4,-1.50316154769E-4,-1.63249845326E-4,-1.75541093365E-4,-1.87171894801E-4,-1.98126221357E-4,-2.08390024582E-4,-2.17951234788E-4,-2.26799754982E-4,-2.3492744991E-4,-2.42328130319E-4,-2.48997532554E-4,-2.54933293648E-4,-2.60134922016E-4,-2.64603763935E-4,-2.68342965946E-4,-2.71357433368E-4,-2.73653785081E-4,-2.75240304773E-4,-2.76126888837E-4,-2.76324991098E-4,-2.75847564599E-4,-2.74709000611E-4,-2.72925065104E-4,-2.70512832876E-4,-2.67490619546E-4,-2.63877911642E-4,-2.59695294983E-4,-2.54964381576E-4,-2.49707735249E-4,-2.43948796229E-4,-2.37711804881E-4,-2.31021724825E-4,-2.23904165635E-4,-2.1638530533E-4,-2.08491812867E-4,-2.00250770834E-4,-1.91689598536E-4,-1.8283597567E-4,-1.73717766784E-4,-1.64362946688E-4,-1.54799527004E-4,-1.45055484021E-4,-1.35158688023E-4,-1.2513683424E-4,-1.1501737558E-4,-1.04827457278E-4,-9.45938535969E-5,-8.43429067189E-5,-7.41004679264E-5,-6.38918412007E-5,-5.37417293322E-5,-4.36741826375E-5,-3.37125503693E-5,-2.38794348944E-5,-1.41966487088E-5,-4.68517434806E-6,4.63487275692E-6,1.3744278437E-5,2.26247609219E-5,3.12589989342E-5,3.96306567229E-5,4.77244060316E-5,5.55259450006E-5,6.3022014014E-5,7.0200408507E-5,7.70499887611E-5,8.35606867176E-5,8.97235098509E-5,9.55305421482E-5,1.0097494225E-4,1.06050938809E-4,1.10753823145E-4,1.15079939246E-4,1.19026671229E-4,1.22592428301E-4,1.25776627354E-4,1.28579673251E-4,1.31002936925E-4,1.33048731378E-4,1.34720285698E-4,1.36021717192E-4,1.36958001758E-4,1.37534942599E-4,1.37759137404E-4,1.37637944116E-4,1.37179445401E-4,1.36392411938E-4,1.35286264666E-4,1.33871036094E-4,1.32157330805E-4,1.30156285279E-4,1.2787952715E-4,1.25339134021E-4,1.22547591964E-4,1.19517753808E-4,1.1626279735E-4,1.12796183583E-4,1.09131615075E-4,1.05282994593E-4,1.0126438408E-4,9.7089964099E-5,9.27739938321E-5,8.83307717371E-5,8.37745969544E-5,7.91197315517E-5,7.43803636921E-5,6.95705718058E-5,6.47042898419E-5,5.97952736713E-5,5.4857068708E-5,4.99029788116E-5,4.49460365274E-5,3.99989747174E-5,3.50741996291E-5,3.01837654462E-5,2.53393503567E-5,2.05522341735E-5,1.58332775328E-5,1.11929026956E-5,6.64107596782E-6,2.18729175344E-6,-2.1594417515E-6,-6.39061522084E-6,-1.04982292173E-5,-1.4474803574E-5,-1.83133851494E-5,-2.20075539692E-5,-2.55514277751E-5,-2.89396650019E-5,-3.21674662109E-5,-3.52305740093E-5,-3.81252714894E-5,-4.08483792261E-5,-4.33972508717E-5,-4.57697673941E-5,-4.7964330002E-5,-4.99798518098E-5,-5.18157482904E-5,-5.34719265734E-5,-5.49487736423E-5,-5.62471434896E-5,-5.73683432897E-5,-5.83141186509E-5,-5.90866380079E-5,-5.96884762194E-5,-6.01225974348E-5,-6.03923372942E-5,-6.05013845288E-5,-6.04537620253E-5,-6.02538074218E-5,-5.99061533E-5,-5.94157070391E-5,-5.87876303958E-5,-5.80273188753E-5,-5.71403809565E-5,-5.61326172323E-5,-5.50099995284E-5,-5.37786500578E-5,-5.24448206717E-5,-5.10148722617E-5,-4.94952543694E-5,-4.78924850557E-5,-4.62131310815E-5,-4.44637884491E-5,-4.26510633501E-5,-4.07815535658E-5,-3.88618303614E-5,-3.68984209147E-5,-3.48977913156E-5,-3.28663301729E-5,-3.0810332859E-5,-2.87359864236E-5,-2.66493552025E-5,-2.45563671463E-5,-2.24628008913E-5,-2.03742735901E-5,-1.82962295197E-5,-1.62339294804E-5,-1.41924409966E-5,-1.21766293272E-5,-1.01911492929E-5,-8.24043792207E-6,-6.32870791796E-6,-4.45994194356E-6,-2.63788772171E-6,-8.66053943434E-7,8.52293023823E-7,2.51413163881E-6,4.11668691268E-6,5.65743137357E-6,7.13408528618E-6,8.54461614496E-6,9.88723746091E-6,1.11604068639E-5,1.23628235441E-5,1.34934250561E-5,1.4551383514E-5,1.55361012017E-5,1.64472056296E-5,1.72845440642E-5,1.80481775635E-5,1.87383745463E-5,1.9355603929E-5,1.99005278608E-5,2.037399409E-5,2.07770279935E-5,2.11108243043E-5,2.1376738567E-5,2.15762783572E-5,2.17110942957E-5,2.17829708912E-5,2.17938172433E-5,2.17456576376E-5,2.16406220655E-5,2.14809366981E-5,2.12689143453E-5,2.10069449294E-5,2.0697486002E-5,2.03430533315E-5,1.99462115893E-5,1.95095651587E-5,1.90357490935E-5,1.8527420248E-5,1.79872486024E-5,1.74179088046E-5,1.68220719474E-5,1.62023976024E-5,1.55615261255E-5,1.49020712518E-5,1.42266129954E-5,1.35376908648E-5,1.28377974104E-5,1.21293721108E-5,1.14147956104E-5,1.06963843144E-5,9.97638534947E-6,9.25697189459E-6,8.54023888662E-6,7.82819910319E-6,7.12277962456E-6,6.42581867484E-6,5.73906284141E-6,5.06416467064E-6,4.40268063655E-6,3.75606947807E-6,3.12569089944E-6,2.51280462732E-6,1.91856981725E-6,1.3440448009E-6,7.9018716518E-7,2.57854152898E-7,-2.52196625692E-7,-7.39306182039E-7,-1.20291285131E-6,-1.64255072004E-6,-2.05784779281E-6,-2.44852391163E-6,-2.81438844241E-6,-3.15533774304E-6,-3.47135242796E-6,-3.76249444454E-6,-4.02890397645E-6,-4.27079618962E-6,-4.48845783642E-6,-4.68224373357E-6,-4.85257312951E-6,-4.99992597666E-6,-5.12483912398E-6,-5.22790244519E-6,-5.30975491746E-6,-5.37108066552E-6,-5.41260498556E-6,-5.43509036295E-6,-5.43933249769E-6,-5.42615635069E-6,-5.39641222386E-6,-5.35097188638E-6,-5.29072475882E-6,-5.21657416674E-6,-5.12943367417E-6,-5.03022350738E-6,-4.91986707837E-6,-4.79928761706E-6,-4.66940492044E-6,-4.53113222638E-6,-4.38537321903E-6,-4.23301917224E-6,-4.07494623652E-6,-3.91201287466E-6,-3.74505745035E-6,-3.57489597332E-6,-3.40232000421E-6,-3.22809472133E-6,-3.05295715119E-6,-2.87761456376E-6,-2.70274303305E-6,-2.5289861627E-6,-2.3569539761E-6,-2.18722196949E-6,-2.02033032645E-6,-1.85678329124E-6,-1.69704869824E-6,-1.54155765411E-6,-1.39070436888E-6,-1.24484613176E-6,-1.10430342711E-6,-9.69360185384E-7,-8.40264164012E-7,-7.17227452294E-7,-6.0042709453E-7,-4.90005825131E-7,-3.86072909296E-7,-2.8870508264E-7,-1.97947582979E-7,-1.13815267335E-7,-3.62938071403E-8,3.46590455053E-8,9.91121276743E-8,1.57159478763E-7" />
// Retrieval info: 	<generic name="coeffScaling" value="auto" />
// Retrieval info: 	<generic name="coeffType" value="int" />
// Retrieval info: 	<generic name="coeffBitWidth" value="8" />
// Retrieval info: 	<generic name="coeffFracBitWidth" value="1" />
// Retrieval info: 	<generic name="outType" value="int" />
// Retrieval info: 	<generic name="outMSBRound" value="sat" />
// Retrieval info: 	<generic name="outMsbBitRem" value="5" />
// Retrieval info: 	<generic name="outLSBRound" value="round" />
// Retrieval info: 	<generic name="outLsbBitRem" value="4" />
// Retrieval info: 	<generic name="bankCount" value="1" />
// Retrieval info: 	<generic name="bankDisplay" value="0" />
// Retrieval info: </instance>
// IPFS_FILES : fir_first.vo
// RELATED_FILES: fir_first.v, dspba_library_package.vhd, dspba_library.vhd, auk_dspip_math_pkg_hpfir.vhd, auk_dspip_lib_pkg_hpfir.vhd, auk_dspip_avalon_streaming_controller_hpfir.vhd, auk_dspip_avalon_streaming_sink_hpfir.vhd, auk_dspip_avalon_streaming_source_hpfir.vhd, auk_dspip_roundsat_hpfir.vhd, altera_avalon_sc_fifo.v, fir_first_0002_rtl.vhd, fir_first_0002_ast.vhd, fir_first_0002.vhd
