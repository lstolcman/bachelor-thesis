// megafunction wizard: %FIR II v15.1%
// GENERATION: XML
// fir_first.v

// Generated using ACDS version 15.1 185

`timescale 1 ps / 1 ps
module fir_first (
		input  wire        clk,              //                     clk.clk
		input  wire        reset_n,          //                     rst.reset_n
		input  wire [15:0] ast_sink_data,    //   avalon_streaming_sink.data
		input  wire        ast_sink_valid,   //                        .valid
		input  wire [1:0]  ast_sink_error,   //                        .error
		output wire [22:0] ast_source_data,  // avalon_streaming_source.data
		output wire        ast_source_valid, //                        .valid
		output wire [1:0]  ast_source_error  //                        .error
	);

	fir_first_0002 fir_first_inst (
		.clk              (clk),              //                     clk.clk
		.reset_n          (reset_n),          //                     rst.reset_n
		.ast_sink_data    (ast_sink_data),    //   avalon_streaming_sink.data
		.ast_sink_valid   (ast_sink_valid),   //                        .valid
		.ast_sink_error   (ast_sink_error),   //                        .error
		.ast_source_data  (ast_source_data),  // avalon_streaming_source.data
		.ast_source_valid (ast_source_valid), //                        .valid
		.ast_source_error (ast_source_error)  //                        .error
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2016 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_fir_compiler_ii" version="15.1" >
// Retrieval info: 	<generic name="filterType" value="decim" />
// Retrieval info: 	<generic name="interpFactor" value="1" />
// Retrieval info: 	<generic name="decimFactor" value="100" />
// Retrieval info: 	<generic name="symmetryMode" value="sym" />
// Retrieval info: 	<generic name="L_bandsFilter" value="1" />
// Retrieval info: 	<generic name="inputChannelNum" value="1" />
// Retrieval info: 	<generic name="clockRate" value="130" />
// Retrieval info: 	<generic name="clockSlack" value="0" />
// Retrieval info: 	<generic name="inputRate" value="130" />
// Retrieval info: 	<generic name="coeffReload" value="false" />
// Retrieval info: 	<generic name="baseAddress" value="0" />
// Retrieval info: 	<generic name="readWriteMode" value="read_write" />
// Retrieval info: 	<generic name="backPressure" value="false" />
// Retrieval info: 	<generic name="deviceFamily" value="Cyclone IV E" />
// Retrieval info: 	<generic name="speedGrade" value="fast" />
// Retrieval info: 	<generic name="delayRAMBlockThreshold" value="20" />
// Retrieval info: 	<generic name="dualMemDistRAMThreshold" value="1280" />
// Retrieval info: 	<generic name="mRAMThreshold" value="1000000" />
// Retrieval info: 	<generic name="hardMultiplierThreshold" value="-1" />
// Retrieval info: 	<generic name="reconfigurable" value="false" />
// Retrieval info: 	<generic name="num_modes" value="2" />
// Retrieval info: 	<generic name="reconfigurable_list" value="0" />
// Retrieval info: 	<generic name="MODE_STRING" value="None Set" />
// Retrieval info: 	<generic name="channelModes" value="0,1,2,3" />
// Retrieval info: 	<generic name="inputType" value="int" />
// Retrieval info: 	<generic name="inputBitWidth" value="16" />
// Retrieval info: 	<generic name="inputFracBitWidth" value="0" />
// Retrieval info: 	<generic name="coeffSetRealValue" value="4.52633279836E-5,-2.78653447929E-19,-5.92639482981E-5,-7.61503615312E-5,-2.19036472124E-5,6.78292668749E-5,1.12924998665E-4,5.85337707317E-5,-6.45569852577E-5,-1.51552746665E-4,-1.10898177766E-4,4.3712519183E-5,1.86027660072E-4,1.77903152061E-4,-9.18284485481E-19,-2.08589583101E-4,-2.55816740965E-4,-7.05454957241E-5,2.10237774785E-4,3.37935235506E-4,1.6959689755E-4,-1.81545233944E-4,-4.14542155815E-4,-2.9560908807E-4,1.13742296652E-4,4.73231413851E-4,4.43047846588E-4,-1.96136053297E-18,-4.99637298275E-4,-6.01898665918E-4,-1.63192596537E-4,4.78575251909E-4,7.57571712748E-4,3.74693046082E-4,-3.95552167125E-4,-8.91296235642E-4,-6.27567678238E-4,2.38557312893E-4,9.81061053258E-4,9.08312507921E-4,-3.41001239965E-18,-0.00100310965905,-0.00119658332624,-3.21377057658E-4,9.33942777168E-4,0.00146555735671,7.18804040385E-4,-7.52722989102E-4,-0.00168300448909,-0.00117621268843,4.43921255568E-4,0.00181308826066,0.00166757771161,-5.18403964305E-18,-0.00181885005475,-0.00215702837581,-5.76102224663E-4,0.001665260495,0.00259983530342,0.00126892869031,-0.00132265676644,-0.002944308956,-0.00204913469139,7.70330994767E-4,0.00313456676138,0.00287297973286,-7.12187138376E-18,-0.00311404219949,-0.00368280684662,-9.81122988495E-4,0.00282952913959,0.00440854724322,0.0021479136046,-0.00223548633921,-0.00497018286442,-0.00345578293049,0.00129827772627,0.00528097856109,0.00484009731342,-9.00131340529E-18,-0.00525116060172,-0.00621654768604,-0.00165844573479,0.00479156309613,0.00748225348859,0.00365534564437,-0.0038165668493,-0.00851710928238,-0.00594747015702,0.00224535851228,0.00918444464737,0.00847082775896,-1.05769527437E-17,-0.00932928457202,-0.0111429182231,-0.00300233533847,0.00877088949564,0.0138664095473,0.0068682775133,-0.00728249373138,-0.0165340451691,-0.0117706387958,0.00454116412054,0.0190344814275,0.0180472137698,-1.16263977579E-17,-0.0212586695721,-0.0264605399197,-0.00747872987474,0.023106340092,0.0390367533073,0.0209430139556,-0.0244921255226,-0.0629093774966,-0.0526159245922,0.0253508739355,0.148707186607,0.261923175995,0.307701100889,0.261923175995,0.148707186607,0.0253508739355,-0.0526159245922,-0.0629093774966,-0.0244921255226,0.0209430139556,0.0390367533073,0.023106340092,-0.00747872987474,-0.0264605399197,-0.0212586695721,-1.16263977579E-17,0.0180472137698,0.0190344814275,0.00454116412054,-0.0117706387958,-0.0165340451691,-0.00728249373138,0.0068682775133,0.0138664095473,0.00877088949564,-0.00300233533847,-0.0111429182231,-0.00932928457202,-1.05769527437E-17,0.00847082775896,0.00918444464737,0.00224535851228,-0.00594747015702,-0.00851710928238,-0.0038165668493,0.00365534564437,0.00748225348859,0.00479156309613,-0.00165844573479,-0.00621654768604,-0.00525116060172,-9.00131340529E-18,0.00484009731342,0.00528097856109,0.00129827772627,-0.00345578293049,-0.00497018286442,-0.00223548633921,0.0021479136046,0.00440854724322,0.00282952913959,-9.81122988495E-4,-0.00368280684662,-0.00311404219949,-7.12187138376E-18,0.00287297973286,0.00313456676138,7.70330994767E-4,-0.00204913469139,-0.002944308956,-0.00132265676644,0.00126892869031,0.00259983530342,0.001665260495,-5.76102224663E-4,-0.00215702837581,-0.00181885005475,-5.18403964305E-18,0.00166757771161,0.00181308826066,4.43921255568E-4,-0.00117621268843,-0.00168300448909,-7.52722989102E-4,7.18804040385E-4,0.00146555735671,9.33942777168E-4,-3.21377057658E-4,-0.00119658332624,-0.00100310965905,-3.41001239965E-18,9.08312507921E-4,9.81061053258E-4,2.38557312893E-4,-6.27567678238E-4,-8.91296235642E-4,-3.95552167125E-4,3.74693046082E-4,7.57571712748E-4,4.78575251909E-4,-1.63192596537E-4,-6.01898665918E-4,-4.99637298275E-4,-1.96136053297E-18,4.43047846588E-4,4.73231413851E-4,1.13742296652E-4,-2.9560908807E-4,-4.14542155815E-4,-1.81545233944E-4,1.6959689755E-4,3.37935235506E-4,2.10237774785E-4,-7.05454957241E-5,-2.55816740965E-4,-2.08589583101E-4,-9.18284485481E-19,1.77903152061E-4,1.86027660072E-4,4.3712519183E-5,-1.10898177766E-4,-1.51552746665E-4,-6.45569852577E-5,5.85337707317E-5,1.12924998665E-4,6.78292668749E-5,-2.19036472124E-5,-7.61503615312E-5,-5.92639482981E-5,-2.78653447929E-19,4.52633279836E-5" />
// Retrieval info: 	<generic name="coeffScaling" value="auto" />
// Retrieval info: 	<generic name="coeffType" value="int" />
// Retrieval info: 	<generic name="coeffBitWidth" value="8" />
// Retrieval info: 	<generic name="coeffFracBitWidth" value="1" />
// Retrieval info: 	<generic name="outType" value="int" />
// Retrieval info: 	<generic name="outMSBRound" value="sat" />
// Retrieval info: 	<generic name="outMsbBitRem" value="5" />
// Retrieval info: 	<generic name="outLSBRound" value="round" />
// Retrieval info: 	<generic name="outLsbBitRem" value="4" />
// Retrieval info: 	<generic name="bankCount" value="1" />
// Retrieval info: 	<generic name="bankDisplay" value="0" />
// Retrieval info: </instance>
// IPFS_FILES : fir_first.vo
// RELATED_FILES: fir_first.v, dspba_library_package.vhd, dspba_library.vhd, auk_dspip_math_pkg_hpfir.vhd, auk_dspip_lib_pkg_hpfir.vhd, auk_dspip_avalon_streaming_controller_hpfir.vhd, auk_dspip_avalon_streaming_sink_hpfir.vhd, auk_dspip_avalon_streaming_source_hpfir.vhd, auk_dspip_roundsat_hpfir.vhd, altera_avalon_sc_fifo.v, fir_first_0002_rtl.vhd, fir_first_0002_ast.vhd, fir_first_0002.vhd
