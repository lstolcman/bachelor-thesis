��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
�쬨����&}GO�X�Դ���}��?VԲH���ǥ���S���8�12h�J�9���BI/�-'�Z��~~�|*z�<�5�E:���t�s�ϙ/m�ha�M��}6_�O`��	��?W�xQ�"~ģQ�M��V��5���B�Pq�Y��O}6�U6};Lo�/1�6b$��Q�wC侢~ރ�%b��q #��q-��C�W)j���o[��c�W�0�A!行���1腡�,D�����_2��ѿLjt0���BTއ��r�<Z}���?���yX9%�1�nS��s�a��+�<���p�:��F9ԐX�]���z��0X;�Â?X��^f��c��勄-(=�/FEJ$���E�@&HO�錱�8K4�H�p1��P�P�� ׼W�C�J2�vV/g f���GO%1�;S�����܄�g6q�,��;��6v!";a���k��J�c$��i��u,��L��~35���b�,f>{ݨ�:w݆Y����C�U�@c����جQWt��ِ{��9�>��-���Cu-!�`	�������,�w��Ԑ5=���k���cBO�*�Iw�Ԏҫ	�_���+�`F#\bbwj���2ր;:$I���V<i�ɲ[�4�f3��>x��y���߃Nh���f-�@���BU��Y���]e���#���\;�	�t�`M�Nc펙fUb�8x�Y3��)�����c6��
&KcQ��a9�S�0�+~�,���؁'�.�L��a�W���J�IQ.��D�l�� �:A���4/B+�ֺ@��[�Mjȹ-��1�Db���BܨH�y1}��8G2���͒$��?�Kp�Y��i��G�˸2謼0��r��o�_t�|��d-�
njEy�Z��qG�s��(6
�W��%�>�UhQINM���0���:�.,��P�B�)���ݬc1�$˱w��1�EdUCv+���}�	I��>�-�+Y`�.�啱��D�)�i���b�̈́>��S���W<��d��V���}���o)]}�y�У�5�a�F��A^��1.3E���1> �H�|+{'����	�z0�K��#&r �dp��j]אtۚ)�҉9�oY`h%��	��x�q�[!d$��0�$x5WY{g����Lkc���E�T��[�����g�A����T�W�>��AG��B�=���(�_���N�8�W� !�0&���Y�9_j(�/_�-Z&D1�'tv�ĥ4'�o��x����Rg�w�ve���h���Y̸��ͺ��K��_l����r�	6������n]�����+[�����N3�M�T;�Y�y?W_�J���"9)Y�KE��^�����)D�2!�@�x��t����H���տ��g�֎	�\��#����T�}�����h40K!�=%����N�vӜvm#���d�Z�)��]'y��5e�+$9�I`B���T�g��>�!;��?`ki2��U���l)WX��?l�]��TY;	i GU�OGfV����x�nU�t���OP7&�v\_�p|'1��	;��J��)��8�a�?��߾�ڵQ����rN��7~��9ք�
.U�]w���X�P?�J.�&�4��M��4Nfhp����Y�[�W�l-���ٵ�]�*(}�n]���4Ch����vȵ���Ԋ����0�+�8�z4O��­=����T����숸r���.�z������/w�}����u	|1�C�����w ���KyH�;��#!��+6��܍£Z)�'X\*%@�f .n	 q�����S��V����#��q�,pU����N�������+Ge�����{3�Ox����-�ji�$���c��� �;T�T_j�D���LZ.ژ���R䝰!�褋^�� Pv�͠7����t-qE6.f4�� YU�& !�
��?��s��<�_B1'a8(������'��ڨr���:7�Q�I+;"u�nY5���s�����Y�zo���rg��x!���DtN���V���t>�(���Y�B��vr�9�U��|?�
���Ƹ��@Тy��{G�
�8�KU6������L�ʠ��v����LopT��&_�`�8�J