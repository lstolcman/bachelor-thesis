��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J�-�4ϼA�IŠ��#�U�(�f���+�p-Hv"�-L��wUoV�5�󷹿1��4��[c��i�>�cű�A<C��'c�|h�H3}&e$zB���*4u����j���YP��
���4Z���UwV5�PƱ�h�u�ҳ�~�0�si��H�d-wt�h��PߴҌ�=
(�@�Ѽ�Ji5�]1���:�A共&bݽ�Q.��=~7�c�
]6�ͤ��G��wn2Ns� �:i6�nm��JB�s���-��#�7q22�}�6sscםy�g 42�H#RRj���3�;{�e�6�]�隬����&򤆘Gj�>"��Jf�}:ʕ����G�,�˙��+��s�E���	KSk�i�.W1Aů����A�hN؏���[_��>:n
���v�6�88|�����_K:�YP̞�7��$Nk�D��ш*�)J��ME��hŰ��:�v��~{��F`]h"���p+<s&�a�C`4y�<%��G$K�o�BXh�Ѯ�M�|T��FEL��/�^�a�Po��K���B����Enrl��t��2�4�5*�y-y����Ǳ�Ӭ�[,�-e�2�����P���~WS��~$�42|��Sw�Y��עs)H��uV_z���c8�:K��|���2�}g�X7H�)g_z��n
���>���r<�2S)��G�(�����S�)��}oU(�*_ݛ��R��ɖd����$ݯHƹ�y���~�*'�d�L���se�
�:#�*A�{��Ψ҆ TΓ=۬=r��:�&��;��	w��H3!y������{hs�H�}�B�!��]Ŗǒ���EO�Q��wch��zI��i��2�%pf���Ȓ�&�7��_��C"�ZMS��ӳZ�&���Ɠ�	�%�
򪓈3���%^0������l�岣�D�i�/��m>x�_�*?�������% ��w�\'�axPjhb��� u�/7� %Uڵ�vu�Zt��|��M�f��հ7�j}�=p'�A�h�MЄ�RT�4�n���9B�6��M�_|˅/�Ƀ/��7\���:����l�RT: m.>� H�} �?�� _'��g��")aׄ�=Ib�9��M�o"z���[|���ԀBޮ>���s�4��`R�P���b�b�?�1�,a�������z$n��E!4F�Y56�?��Y�+,�JӋag0������h8�B.��_j1C��܍�����X�U%n,i�ӵ�
��7t������r�oF�$����B�5IsO r�J�S$��*��Լ=?��RG��Fv�(嶱� Y��lG2e��3]��4��/�E�I�۳���l�bQ���o�E�����]�����.��'ja"�u �� ��}Pn2�Y��
n��uK���JhO�� Ö�}�$6�`K�WI�J��� կ0����$��Gwܵ�+��	ʽ�X��n3?56`�)��w]i���B1�,���pT�#K�%.�~r�����e��E�/�@bd~�^��d�ɞ���b8)�i�PBc>qřگ3���т���ƺ���c�̃��H�A�ȹ)OY�lκj𚨌#��)�5��V�צo#;[:�TKk|�����P� �R�Z:�����nU�����؉!������CL�1���$�i�n�a��C`	^Zmb&v^O����nӘ��Յ���D�U��n
��qx�.T���nk''nV���=��j�%�E����6T�{\�����us����Cf���y�W1��m8=����qĜ�� |Mrȼ�H��}��}�$������dC����iA�����qo�d�KC�v"YSQ*��4L��Qq�������!N��g��B�9�3+i3A:|ږZ=����-���䚂����펿��s$����p�p���������B��Q�o�K�˳��X3�����/+�M��C�*��Ѝ���|�
��Ѣڨ�^6P3;p,@��y� �O�0ȓ
Ry]:�N!�+�c�������cH"��F�69��ۤ�A��b�>�
�O�k�I>6�ޟ �(���-i�A��6����_�S�^�U�B=�+u.�P����� xDɪ"�G gy���U�!�^�CxٱfنO��lсZ���[���['�,�:��2�lю�qt{M31�6Sd��	�J��.��@�Jatu�����G�h_b�
�* �،�4G�<��`��׷�>�R Y0�����xR��L���i-�4[.bIb�ǧ��b��s^�F�T�-%��M~B+�����-�O���,��!d�y�
��'����q,�����G��ڗ���T�:O�p�P�;N�{�8�f%�{����@uI7����;N�s�M�R�ط�{�Φ���Ͱ?��T�y9�%�W���o&�����F�yv�3���{{7���K��n�zN�j�r�c��/u� �L����O'�W( žD7��_Ԁ��ub�����S��v��3��e.���xj�8ʇ��왹�<������Yi��g�9��*��Ln0�1�q�=���'$���w-9��S����=��P��k��`��Y�\j+ ��*�o�*,�*�7��A=��Q�_�\mAX+o�63��h��=�P�<�������p��ق9����+,�HxQMn����6��N%W� ��i���t2�c_�M(���,�K.�C[����K��p8�
&&%�C��X`��C� ZP�b��o��ڡbͳE�uz&�)�Z�H�ӡ������M��`ԚZA9���9)kղIg��ˌ@&�N��Le��'׮T�H Q[pQub��,>F�d�#����������'[�'j��⾈�"�<؜��NNU;>L�i˞�R&�"���S��I�ź��=��ry���O&U#��-�Ac�n��⺚��I�l'���M�M} h;p��8x��ߞD�<2u�Jw�>����Q�]@��¢�ࢆ���`������oS5J';ßw+��9�1���[�} �����|��Eg'��83)��0�[iM#b�b���<X����M��݌��r;.��z����m|v��Fu����Y��V(�Fw��vh<�ddX~�wf0>Nr�X���ʟIH�;"��V�7��0����N��U˻,�L���\�c0S������#�}0����m���e:�)��xW��쌗���J&㞈�}�'d0�q��%B�w�>P��t2% �`�P�4�>���𩗠���wN;>����l��`�R��� ����9��(��W$:Ck�g3�W�Q���d}�hߔ�S\`,���/kt��|矹���&;���%یR�`#�'%�B���LEm*|��r.�y��9�Ur���A�E��q�����g����;����@|?4gy��:�$�]�~=%윇�jX�]�>��r�Vx�C3���{hh<�L���>A2Q$�JH7��,�r�6Bv
����]e_��F����]�v����2��^/D�n�vC@�[�!�N���,}��v��s�N���D�<�8�� ���K�X�#�?��;mܭ�,��S��� U(c��8a�*O��L�$V!���8�y���"�e�z_����.coiy$ }�}���%t�Ȱ��i�I{U�un���9ޭ� b�Ċ��W{Z�c�/A߰/�Q�u�?�ą���	�΋�ȋ*G|.@���Z.e~��94.0?,��{�w�ٖ���j��ԑl�ee���%��7���,P]��AR4d���
�ܽ��hk���nx/Y�oYIVO
re��Q�	��� <�(�@)�O���vcgR�� ��0/ ��xBx���Bۤ:�d!<�J�R�W3-����a�B�&���G�M[PF�i�6+��e��&�/98T��_F�ːVopm�������䪈���6v�ӝQ\`�m@)�QBg"e���HM�*�t!����?DS���#т'�o��!7Qa3�BS����B���jg�;�<$�r�*��@���o�!Z���+=���0�+�=��W�e^O��pt6k*�Nc�.��n�q��"��c"	���(|�e�E���:x?�յk2�qGa.|�˥l�h��d4_|�G����z(��vmv����f�,h�G�7�����[��w���0�Mӛ���]�=3ꕽ��M/�>����,Q	k�OZ$|B'��?�m����ț��35.:�8ZkԬ�\�?��u���(t���*?b�~ޓ�A��m��w+EG9���h�x*-*�_K��~���'6�}��F�M�C����i���b��X���M	��y�Ȃ�=P��@��K~k��l_Q�p��i!7�Ђ�"�<d��S�9��Y� �Վ��S���D�+:�i���bP�����VΛh��k�ME�,�U��PUoL0ѝ���GX��蝋�}ك�. u\�����6��Aq�%�u�a��$�^���93}�.F-�k��c٦(��wDt	˟��}��cwƧ{�(IA|�`��V��shx�����.���E��TuJ�!$o�E=>P�rb|N����gXf�̈́��ʰ����M�/���DQ��>��E��`;ވ�Uεy0I]�-���MW��^�Hj�^��Bܞ�t��|��_�'���W@w�݅�D]�=�`p��tN�`f��� ���e �o��X�o�ֆ9_���Z \�e*�mo6N�:��g�|-+�P��j�[uX$5Ӂ�t�j������ �A7ؤ���!�K�T�	Nd~ҾH]4���_X��-���sV�L-ث�G^ִ�I��M��5�4�NZ@�"N]+�5�o_�(fH_�߽��������ޒ��J�[ �8G��B�����)��ȉM˂*��uQ��b�آu�_�uR�ǏS/h9�Ӽ�;F�tz�T�2��|a���s/X�9��(�wl1x=p�_۷9�y�3�:���8F�"�M�_a��6Ѓg����mB�S���@:�|Q�rFՋ�w�VU��hιN��,(���8Ļkx�2}�襐?B��m��aC����eE����.�=�3�7�L�`vY�����N��/:�N�|�� ��K`ZU~h��A�yʐc�dPz��+�J�/�v���K�d��e��ڄ���[8Lju#���6�	���8]��P:b��ΏA�N��	�2-�,�^ w+mR���2�ܔ)ˬ�Ի#�H����U�F6-�0A	�����5�l��W��	�e���5��[�z���6R���n5)OY�o�6qǹ�w�,F�,�'s
GL �/���1��p3/o��K)s�T4.��5jƍ��u��[��T�g��,P�3Mq����턷 Y犪;��h�[x�5w�`�f��a+�����X-���I��Z�4�^Cޖ���ԛC1��Po�k]�ÀJ�����{�Z)�䈌��
l�c--���l��2���� �*�0�wdo)0�{-|!�M�J9�\��l�}��*4ad��ߣ����G�%��s��|��f��E��}9�>F��� ��f\�\9�SE�8���b�1����j$�`F�6�ͩ�L������OZ)k�4F�����Q��R�h8[o��C�
�"Z� ��z1m�Ġ<��d�y��jyC�}e�a�,N.�|$k����;��)�/�~��E�E�~���A�z��~df���C(5�l���(��덅�	@ޤ��Ho��5�Fe��<���@P�6̐g粕����ck�1��=�i��+Q�*�x��̰,n ���"�H�1�*����y�WW#�n�bPA�a`:�vS�B�F]��c��`u��4�ڂla���f���c�4fR윔m����|�W��j�6�f�Y~1*�!ፄ=�Vۼ�X��ߋ��]�~�F��G�P��|��Ze�	x��4%�z���5s���d��W3��4�cU�F�)A����3��c G�Z��aM+������gW4?dy����*t�,�<�tw:�~��1�1!NU���?����3��Nm�x��6��PsEf0ަ�$���j_���ˁ�hYh��,g&I��}�;��L�S�4AI XUa̩]
�_1�1�룁d>f ק�4kĦu��
�-^�$-����uC$Ͻ�>5$�����d��~X:&�]a~���5}^È4|�]<A���F�(�������f�*��Bs���l���P1X�������X7N�Xjە<��y�Idq8!�q��S��KX��I�JUEp��$o�e�Fܲ��^�� Х�Sx߾��Lƛx+�<����H��Ϟ0\`-
.~��C�SJ$}(����qM98	�H,K�0�R�M�t���5@|p���$�቉��pWѣ�I��A4��3�X��y��)������]:-�܎�Y6�\��Ik˝j+����oZ��Ю>�@�޼��y|F��?��I��l*�+fd�x[�;+�׾R�S�B��>N�ʌ��y"E;�s�ؐ�����#/pH�B�Ih@#5�����3�	��1=|zc��>|;*�%�ZV&Ż�l0#v��%��G�BuA&����]B�Z����`9�)��9F]���-����fr�;��H�J�Mԗ�P���.�m��WAU]��(��$+P]K���۾<2��(�#���f�"�f}��}I0舾*x|�����Oȉ7�E�\;~Ө����W)�x�j�4���1�L��c���}(��R�5�����F�d�:R����\k�+�������a�Ǣ��F���]�wꏨ#���@!��x\l ���5s��G��;�p�'��3����p�6��:�$�	�z�d/�M�P���wj�ۈ��d`���2p����,&�2�*����q���`P�%_��X-�O~_㘜��i݊1��j"K�\ʫ��F���x� ��qW�=�������.��ť7w�S1�y��m��Sg�)�<]p�`0�WRnw�tA���i��\N��s��n\�� �:&[O:�#ݵ=��A0�o*S2x����=�xU��� v�kK0p�y&�V��EBO�.~k�T�p<��q�yo&����Ry�풫[}����ZF�L~Q��m������ҕ�����q������N�Gzc�ƹB<���M\�mkH��3�Λ�&��WD87�杍y�e�$��v�R{�W�\
��~�ٮoG�������Ks$EEC�s�q��ٗh|<����<ﮣp��D�v���9�ⶏ�,�G���3�/M�eI�"Gd�1t dX�
�H���`x���㩈�i������~�xw D����h%i�X"!�~��y�Dx��I��ձ��y�Z��Od�[do��ܴ�j~s�nFn�l�9��L���U����3�k9�/)�6FBU/k���N��XJ+Y