��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J7���zZ�3������B��h�Y!,�c�k&^Pk�����[N�w����$���/�bW�/����F�@��=�\T����&#%�,:b��B���K���[��BzE���|������B���ʫD������X���^,J����xGO�׾~|2����/�������n�3���r��]C}��miA��@�\��|>��pZb��THx�y��+��=����߅.��Ӕ/�f��E�3M�����jX�H�'U.FT� ���J�~�.�h�A�Pј����'n��w���.솂nm��k�6�t��性��+煠�D�:�&��5�X-���O�u��r�@�D4H'�O a.��B��Ty�b{g��mV��d="��y� �;B�P
`�,_H- �Y�ۑ�q| JZS�2�!˳S��Hꅙy_�T��!Y�*�V�\w3F��[��A'������%Ԣ���KNK^}�sV�U	H�:�6�{Try냓�oNa%���ȥ�%=Rx�A�q� �$�&�80���h�j���-qv�QV�Ӣ�\$M��Н�k���A����������ze�-˘��j ���������o��M{�e��0@�$�v���8T������^5�4��Mi4�[
�`�U�~�߇ �I����Ɓs�b�2�),����s8�]��+ci�e��]l�����So�������D����{(}러:u�޾=$3�d�\��͝x����+xo�O@��B4�RT�,��얔�F�����6F?_�/}�	1����o�q^4R�`2�3�4q�	���(|Pwb��Q���;�Du9�p�m��qC����M���K�R4�1��/��Ê<?�l� z�cm R��}�D	}=3�lJ�9O2r�<Ab:�GbT_i��$�v#=�/�U����9y��v�MۂBP��si�O�"�@�������[������&݊�E��B�-g�/y�e� �rs��~3f40��{\��J�1"��Y�N�_�	�[�5����{%�k��Kh P]��/+?�@p�(�I��Q�ظK�c}�������� �u��;^8!TN	�C&�Z�M��ځ����O+U�`���:YF���nLW�`M�){L��?�(d,n��Ġ\�5���$�/���A٭��)�o����=� ����R�0*��.�M���U+��s�jl��hA��
�i�P����0�Zf$�]��z���G{��9�T?�>6N���%��Mi�F�Lg=���tl�ȶ��-�
."(Q
ZY�ɉ�O�v�P���F�U~��J;s�h5(�F��A�L�f6m2�����y��8�7t ��7=�AM(���W�4t
��ו�p*�߄)iY�S��nL���~�q��~Ď��6�ǽ(�~�"�{<�<9��c�B:&��D��J_]ꑘ� �W�ʶ�J����X}�DI�e4�:� Ado�UI�!h�h-�e-S���k�V�k��ot�����F5�+C�ڄ��s�H	�v����#s�{����l�q���߮P^���X���e�~�����6)�
�Kڸ7�VtP���q����H�ˇ�W�������5Ʊ��YOLm����怽Uƶ��E�F}�
�������GlZ��Ly�����n�y�->D;��W���������E8���X���d�7n� j% �C���3���� ��ݛO0C{�b��ދ~��Z�fq?�*"_s���LT�彩��~�b$q.��d����$9�D��vO�X��v��~yS���� �h4��V�v����p�0������,Tj�;��tU����F��ka,������$��-֒��?����]X8j!�˞�6_���BI���`�Bb��Q�n &�S�uOYD���NS�)��5�I#�=mD�r��q�
z{{(Y�}���[�h�/`��7B!9�6��A �S߫�I�Q�a��K$UDSۢ�:�+K�2PPn@�K��1���.�� o8?oZ5/mX�\��+e�w�5[��<f�jc�T�Y2l���u�&hegPG	�A-7�8e3o=ő�@'�_����!���~�1��,�^b���mϼ�|:4~&����*��s"���1����v�Xom��r��j!�x��W�4���DqAe��yS�I֊J^��ꂈ(�cs$�JJ��3��z�3��>����Ĳ�"�s D1�p�)=l�FB;�8Q�Y���3׌/�r�;�MIh܈J
8^�_�D'd[Ղ�t_��W�=�-b#�A]~[V}��#b�>���dp�
��+(-7��l��X�:P�AȓзF��_Lt»����8�QL �6'��^�D��a�i��?D�}�%����I"s�'�g��߁/�0x1���_��:`Z^Ve��SP�,���m��� $�檲0��z	�Љ�Y.�t-�N���X��`���<��O��N�q|!�}�`��A2=8:	O��t�e-]�z����'4�3̑Gobl�n�P�~(���S��Vkt�p�Wב���~�;�@�!�aĚc$,y�0���1�{�����`J��/kBzS�[s=j������]�Zv��)G�%�ۥ X�;���zI�H�0C��p����VS��[Cy��'�X�����kz�_���O��듑���iS�Lq=x�x>�rx[�����:����ϗ��	�Ze���xH9c���=8��6I>�"s.&�2������Y��S�D~���C*e�q�Z��ĈƗ�[�2Kܯm��aH8�zdvIF�-p3��[�d��y��;@����Ц�@��i�YTc��\�s�T7
��F�?�2�Ǘ͠�N�
��uK;
�~�(E���7cK��>��7-�䠃�ڀ�]��k.`<��s�_=��nZ
�d@�&���4���}�~�e�N�#���E�m��ɸc{�hK�/���!����0�r�~��§i^�\p�1��o-�Y ���l"�=1����ޕ��g-s<�2f��뵳|	M]cQ��Ip������2�fH���TU�}v��	 7��λ� ����aÐ&��ې��!��[�t�s�_��Dy>w�.P��Ro��@E1�ߴLU�r��k�+wO�_�WL}F�!�A�O��i����_։@1&U��X#�E�6ja���<����g]z�I2x먵r�6n[wj�ӏ«=�	��Ѻ����*3]F��QX}#6��}[5lחЮR�q~R�z�.gF���M,}���#����3��%R�6U��M�R�c!�ms��[o��}�b<&[p˷���r�{�����<�fi��%�WK���iث�򢅁�m4�(	�o���Dĳ�*T_���Dk5$p�xsR����b�x����R�u��j��Oh1����06��e�%��41�|N<p ��\�ٰ����KC�u8���^�"h	�;��r�px\����B�U�_Ey}��oݼ&�#W ���9�5�����(ʫ�[qE��KT��T5� �h�h���|o�*^c3՟�\.2�m.^�#�]��:ھ^Kq�7�:��3`���62G��i�Ӗ����s/M���m�=�x�2�?^+N�9�~�Ȣ��S�|3\�ӹ��d)%��j<��s�$@3RM������IM���0R	Ɛ����W׋��j�*�������s�+��1)S/�O�I��h�ݮ�oN�1����F9�.F3�6"(��XL�o�{^���Ӌmr�0�J5��h�)���>?�o�� �4&O�����^�%S��07݂�8,���0�$����EI���)|�\���Ka�Csص�����0H0�t����P�������.�R���c��E��-�� 䕂	�:�Y�JG�'��9GpUo��\ ����#��!�ɟ��ʙ�!Ge���҅��Z��W��a��E���dӕ-����n\� ةG�r+���Z\����K�̉��Y;�F��՛US�u��	�R` cv*:�Kق��>Zc��v�>N�\va n�;�<S2�aA�u�q�[T����"�D���C�	��B��S~b�� �F��$�dٻ?X�٘eԍ1m�ө�L_U�v����Z���t&Uʵ0�����dz�T˯aVA�_
̒Q����bh���?�2��A��Y5~�-W�Th����GՀk��kD��az�c�WfR�y���gH��O���5�0��q�Ͷ�py�%3�"�|le��k�y&�σK����#k�B�$d^CV���ϦfǱ���ܺ�g	T��.�S:k��I�����G��s7�zfg�ɇ��6=R�()�Bԙ4~$+b�U