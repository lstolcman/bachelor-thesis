��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�O�5t�"�/�V#�bnQE{C��P�oHȥ��S㌰��'�@���:K���J�7&V�T����F]X�J�ʨ(��̰͑ާ���bރU����B/,d�{X�F_�@�v�k�7S�x1�=�2�T�ޡC�� 9$<3�W0Q���a�.+:��JK&&N��*b�"�X��)��+�t�a���:�	��L�{�V\ث{l�I�����T��d�l�o��ir�4 $�X����j�k��1��� �?������%ڠ��3x�.9~���e��S�*�0��%2������eFy���Ż�A7W�`'pB�����gO02mjV/*��ed S[�Wk�"�F�e]�O��V��u�GzR��7��.L
(B���r7F� ��ǽƈ��<i�SE4���َ�>���I�{�s�3uQ�j-Et����߁�Jt�OoV4����Vy�cx���5��5�|>��աc��B:���|ƃ�v{5��gg��(��S�� }E��힒��p}}:��_�{� �):NK߸@}J��Gd�T=�y6j�ݯ�D���
Ƹ�����{�H1=)o��AkRZ=Ug��&�%��w�`7�%��nd��@"v�4�w�%��m�	��g��%�ӊ��:��
%p��`2{J�R�I�9�Qt?��4�n{���hw̒�r��K�����eQޔ~�l��/�C(HH��ĉ��H��������u�%�jͨ����s�ޱ~���|Cq���L��qϤ�Qmb�+�SAh��;�η5�ڱ�=�j�'�DM8O6o;�x��vK+�`�u4��������P9�_͘�����#)F��	��?m���Z[2�I5"y�K[�{�Y��B�7g!��N���&���0�g����0���M�=UBoW�ϡ��W0}�Q�����h��­�7���{�ڶ�{k��*��C'����׾y87ψ���ޫm��rQ	���O.�]}Z��Y����Їt��.���!�Rѵd8s�^<^��6u5��ʙF��Vݻ��*������&���O���+�q\K9;P��ə��]���POM�Ϡ#%��k�I	
 �v��p�{{x�_X�s�h��A��r��R�RCq��Uj����D��۲4(�W's�w��g��	��3қ-�:8���r��H'.��#)�G��t%R�{)쪹��m�Q�Cx�ߩ4�4���ː�W���s��~�z㷞�>�#�}�i~���C8���/�/n3a9���US��1��nv��yj���
�ܥ�U�,��6���U������V��P�� ��Y�tW���&�������ա��͜S.	 zm�a?;�sk�3������l�3��n���*ݚ������5�Z>��΍��9�J��.��ir߃�Y��.-�5G�e���H�; ��h��>M�;2,���V����i��iHh�*��쉙&Г#R�v��y����T���K��&���%��0�hbˤ��{:�C��(�x��tX'xl�ZY'n=�o!
�;��6�#+MP��j�(Y�a��
$�G�����!�m�j��}2���C��0������[փ�)xs]�aKj�[JW�YJ�ǧ�_5�qrr��/�&&�K�[[��Y��H���ŵ�w�oF/`R
ې"YQ��Z�*\#`��� ��J�ΩԨNa`�ߤ/ʦ^2*�_����x$���� �m�O��<�������� r^���Ϛ+�*� g������ؗ���@|1l���8L�V���,�i�ƀxz*ZȦ��k�I�̐W���̺�8pl|gIs�E�b�kl����w����^�{H��A���ߥ���xT3��l�PV��B���)L���I�	��#_��Iq"�:ݏ�AL� ��U�]/�Q�����w2�.G���XQ�ጄ�d,�bΣ��P��?"���߾+$�������A�n/���&"e�PlH�4r���? ����0���}���*��纥����|�1�|f)����k��]WO&X:���HH�+�O@˵��}Ґ�fI��� "���뜋f^�_Z��a(O��p6e��`��#�������vN �6��Iq��g����r��������ٔ�ͬ����,�d9�)�wxc��,�ڞ:��MP�`�}�̈*KA�o�ȆR�X���^����"4+�4$;��ׅUߠ�"yd��%NQ�w
/�zr�4q�w��,�eY���lj��1ά\=�om��ZѓFV�B��k�|sc������g�6��O8#1��2U|�6��� j���g~�"�i +��&
�ϫ��-F�J�Dn5Xh�Խ��1a�����rΒs.M}���wa��� ��c�� 1;�o���%Q2���,%�S\z����b=0�4s.����J9yp2�;�,m>�����"�����(��7D_�0��B ?��7��(�ռw�4v����.�	1pO41���,9�t���3�b�}��(Y2��޼c�*#
�^p���\�gbn�'��lKr5����8G�I.�����"o� E<�'�b���~*(�ۜ���L��K|65g����t��ƅp`����*�<47'yܵ�o�]6�D�ɖ`F�	�@}�/�)ȼ�X��ld�jK9�������&!$g��Ǭ�.B�*��?�[F�̪4�ā1�7��l�h���r�M-F�٭��U9&,JY�:�7a2�L�/6T��*n~>'E����h8�3��쥎�����1�\�o:�}K3l�j/߁w����^<?�+�s@x3ݭ��jЪ��y���鬫�F0�$R� `gI�͊$V]
O��Cn�}:P�L�K^���y�؎1*���嗐I�cz0`���vo}���qZ^0>8�2�X_���Ǉ��b��c�F��*�yC_0X>�mz>�Њ'��Px���!<�F:���Pv`AN��W����v�Vm���M���8��9
3	@� u#i+j+l���j�J�IFᡳvCM�����:�^ua�;]�q��2'�n�+�%�{sܺ+��NZ#h�&�z�uQb՞�.��?q�o�!�>��\k��C�.鷛֓[?�����f����>Y�[9�!C��e���B���#_�ц�+c�t���o�$��_���Ŵ>/8H�a ��.����,CN�>�dT��Y��6��x4 �}b�:rq&�5�K�N�f̿�U�����|h&a��u?���8�k��UC��Ho���s60Ry�U�>��v���n̏��?�nz���vq���(ڵ�Y�8��o��@}h��h�\^�J�d��#����ư����v�[�7�i����� ��]�0`��l}��j�a���U��"����
b_�eWB,�.q>S��Ls��ň�MNM�ݜ!rE��02غF���=�������M�����|�4LFd�11�F�ۣ$
]J�`y��y�}wڠ�)c��LB�!9��E�@��yGѱ���!�ٲM�´;�
��
���)?`�|�oLyu�����v��`�2�R�q�7k4΄�KN(`x���q<�P.��}���8Ӄ*�T E����w�eyL��x��ǹ2���!�-b���Fn��f�N�p�Õ�l�RO�g���&ZD9ۂe�]]/�A�}J���Z,��da=��x�-!:D�޺6ono%����/�u�,-�v�B�
-fQַ}�d��@#�4Z��R��:�%]z���]��	��+w�#pKU�n��IU���q(^��f��:���qC	4�M� ��{�F$�v��lH�Aܻo۳泸���'�բ���g�4Sʺ�l���A�����$��|L&vN$A�|]�Pv��[b)wz���pK��^)=��B ���I����n<�r�*	~^��%�1�Aq�c ��O�P����j\XlU�hV��d�Zs�p�6���Kۣ�����9uk�DB%��5C�C��	�<�����jl/ږ��d{8gv���$~�'����1RI�5uIvUG�}�fnn4�x��� ��Rr����x���:�.HT�����E��w�tP9υNK:v�B�����]KR���+�M+r@T����r�-�W�r���"0�Qݿ�����oJLwS1���d�D�j&�F3M4\�yWg۫�6���������B����Ts �Vr�4�����mfZY1���j�$\���ҝkC���D�3D���|�d��
�(�>�X��'1��6MҎ �����Og�5�2�'��E R��,�����=c����bn��f�)Z`j�&M����xb���>o������M6M������.�����v����y�*ϑ�wJ8��o��z�n���춮���ï�V#9���<�pЅҍ<�����!�Z���oI�°$��fն̙&=K�|�CnfL���!�q��.£CX����F8�9�2�ܷ���,��9��^E�8eIe��D���
�M�杂���?�/}K4���
��$M����}�l/ N�#SJ¬���q�^ w!� �Aa
m��Voח�Ǝ>�ŕկ&�T^�<(�&��m�a�+�&*�s�AY��2nufsF���>W�?����5�5�o�_`�Rv�90�6����/)�Uя`�F�,w0!+��������E�aa��!�=��Wpl��Krm���)�ᇧx?'�E[�"���5'f����B�n��!�D9N�"���'Wj=6q����g]�0��+
����B~]��X��M!vRK���s�c��:�0TIs��6׾�T���$o8�֨"�����J󶾀�A�]_W��������77�.=��U�,�'��^�Q��
y�Al} M��cO|̦�_�qjB'Ry�H`�`
c~�˖r�'�v�?�$�3�{�1uQ~c��D�8I��^�|^���XIt)�t�6	��?�¸�*����'!��
dT���,_��ԄՁ��^ /���̝N�Yʭ?�~ٯ2X��i3k�匾�V<?�ČT������R<�.C�h�y�[\P�߇�-��W]�� 	��`&���_��ߚ0��t���H�k�,��@u���a)ѽXe6�)�mz�U�Cg�eVa,�e������fI�σ�1p �=�2m�)q ��<�ؘ��̘ˠ�K���!��Ȕ�v�J��Gk
�N� �ٱ&�:�1M˳̓�m��`F�	�dF��v���Y��"�	Ws���p�Mn	�b�,�wM�!���I2�3������@U��.'�-�tYj��oD`$���ѭk�֔$���I1H(POBe�a�9{J�['�i��<8��no����y�씉��R��06Ftf���8'}��L-^�!�%�"~��6�u�9�9l�!�����n#ZY'y�M��j+�ӆ�|tH_�!,����=n���{�Iυ'���6�@�ga �Ȟk؉��E�Ā�5����jt��'�K�H��n���֬�f6L�ud�+��.y��cKzgϰ?�����6�O-V�����Lk;��-�SU,�f���������%�\V�N�����s�N���m�S���sg�}�ޚ��*�����n��. j(�z8O�wv��\rq4_�L�j�?"		{3F0s� '�+q�o���!ć����ky7]���JGg?�;�8�����%<�3���naRJT����2�;y�.P��G�֎x9Mσ�B��w�o1�=����Au���e_6|u�[X@`����>��1�f��8�d�dseW��C7/����,��<�sO���`+��e���g]Ke��q\c�&����4{DP.-������b[�7�h��_��J�C�^=�d�~���ש�R2����c��.,^И��5��F�L_�3��c��&���s����Ͳ_x�W] 6N�p�u��i���N�"���}]��_]��z�*|�n�����$L;�a~��a	эU�����O��>u}h����8"�X�T�Q����)#7�Z�֜/�R����"��
�X����k��aM����{�)D�ƒ1����J�[��8��m��@/����Ix'�>~�ko;�����]�s�ba��#Lӈ�J��S�"9��
_�s6y[I�q\�+a�����EfYo�e/�'u�v����5�5���1���J���O��.pv"G���0_*�9�~�T��<RTcΜ���G���4j� ��F��T��s��Z��a?)WGv�,��A	eM1>xd@�R��۹^=��\���w´��]Cm�����p�rY�����'B��>��Ix{7��B~3:����]�G2;O��%�IL���r|�<��P���A>��m={�g���~��`p��Ʈ]��'B�9��a��p�'C�|�#D���cR�	J��t�'�.WCvǹz��a�9'0t��a�)��E,'@����+}GPȊU$JR���g�@��Օ
4�� ��~��>�_J<?9�l��"ҽZd�c_���};���N�)`���{\ø-�b��
��Fҩ�w�����q509�c��v����c�}�T3��9%�wa�!짼^Q�v���k�[�@�8�rj�� �U���E�m�u6�n�Υ�w��R��m���1�Rङ���Ǭ�{!:Mg�T�r�O��������x��4=���I�񉜴~��$��a����}�����N>�[a��s�������� _uV&����T���R���D��$��RA�b���U�[�z�J����t��[�gX|ݨ��8�4�`eN\ݠ����E9�AԜ^�7-߁��ط��k3E��P�MO2#ʊi��]�0�a�^p�����N�~ @;!��J��rV�EP��5��������˰@��e� P�qzg7�Ͱ��h��L�3���1>
�����n@� wmp�
J;JOR�?��t.gA��p�<:5x�γ��?����k��hc��c���i���,8y3�7�b��iPb����J�V��.�%@ǰ8Hyu��ވ���օ��/�&Rc��۽���;H- �j�PB���e���Gk�	e���k��@2B�O�����޳�e�ОSx[~�����vo��"���.���{��7*�z��z���E��j��d�|�$D��\����e�26�&�'�ʬ�a��\��r�%��)���Ml"	��z���\�^�V��W�7	��Zf0��ҥ��Qal��,����i�uk�-fbH���F��8T�GA�`s���|����*�/�T?�CSU���ĸ��O��)���w�]4w��%ء1Z%ǁ��o]&�G�Ӝ� O�s�g�����۝�ھp��=���%s�͓������,¿�*��*��#�CRy�$č��?y�Q��s?N�#����F�_��)���JEe?^&���q�ο7M��zգ\�]6�ۿ�摒N�bt��G��^�����@�jg�b�y|h6O����"�0���Պ嘧zNK~]ŵ}����V�fϒ(:��G]q"WB9��5������*���2�[>f�e�xv15	��,v���[��)]��N��~`���z�뷨P2G����+h��.]^-6�� L0�p\�B��ipr!N�# !t��C��������d��-_%p�U��1'>��3�!x���z�#�QA�eC1�㋯�}��3Ih�&C�]{��.�d�]ޒ@u��uո�����p����Uˋҁ�%⪟�5���D�l��u���lȋJ0�h����W�[t)]�@a�K�m��⢏;�Kno-���v��������/��ˋ��Cq�@��H�=Q����^*�^ݩ��ً�<x�c_���<+�a��uaϑ̔��!�P��\��<�)e�Rs頚�VҨǙ�܎|"xS�J쭘�.���k��Qr���S�ĽH�Ex{��ԋ�b����,�È5�M�0�7�Mh��a�5��ũAz�'L3��rZ�OH)%�yc}�%�5���^�d�T���{�-�ܶ���Ћy�ӏ��G:u �$�cKn̊���QD��?����A1.K襬K='��
�U{-��7OW9�\�-�!��i�D��GTu�*�]�:���W���Z�CVi�g�Us|��T��@*b��5�����̨��#�n�K�*��B�LXM�q�1��Ie�RO�շ{��,v�����#�@�UگuG{��u��M.{c8/T[�<G�"�
�`K:�~�p���\��6��ڗO�ƙ��n9a������Z�lt84�UV�L7�����
5���:��*�$���hx�Oi\K_*؋��&��X�M�S�A���v���Bf!R:N�I�}��^����#L{�\���Q�ws5�{(��)��7�=k?��0�G���ƻ�g���&�f�>�j
�\�x��ŗ�O3s�+�M�Z+1.� խ�Cf����P_H2�e�5(�q�XT-��皏��ى�ʓ��*���)��4����~x��@m��Ū������^o:��odPց��;P��Li�1���U���U�j�v��	�5U����I��y������Ȗ�HNi�����Qoқ�X�D�M��192�;AJ�����-~%��˖i�K�<*]rɑR�*���p�pZb�{е#"r'(���vV>K˦LvY㗝4sp�'�:�o�V��.y��Wu����q�6�o�.E�4�^�}��Y�j�rN���Z UVgNȈ�^A�H|".|+���E(�����T���Ŕ��!k��J�>��V4=2kvR2��q���!��}�~46�%{̶��Fn�3`B?(�$�I#��p��=␎q`̀S��<�� ��za��Y��vćrY�6�Z��˂d�R~uG�o��ؑg�WAV<�z@g��k����"�U]1Y5ʯ@��D��֜�b�p�ԑ�?�5���CΒ��[����`����F2w�V�L���i�F���,T�X��i�p�)��\f˩�?_>�kKe[�0�$|@���y ߑ�`JJ�VO�P�:���Fkw�3��'�o�wi�4Q8:	�.:?��2�6�ِn?�����(�'��o�	^�!�C;{�YЬ�����Z5O���_u鞝�޾����+�;�+�:�y i�Nw�ڻ�Y��-E��|R)�c�����!;Ұ�Q��B�OoL�f�@@���ν� �^�4��ΓT��\�����ӭ�Ĳ�����,�-%(�0Z_�H4_����4��xk��֮ U"�_���H�|xT�h��M�+ %�>�8\�H$�T�a�bMu&���(b6�����]b�ϱ8̾��F�]Ix�5��-Љ��Ҟ�l�r �x���]�@G�ׁ�I/Ū�8� ���V��3E����X1١ɵ)�őUP���1�60�d�'��ܬ�C���ok��`tjy]����wd1�VÄ��L+����Cq�"u��؀����uR�q�y�}x�iԽ��諊��ܷ�9Z�����5��x�_��^Qe3RӶ-�.`4F0�
���^A�F%up���N���㌵���t��բ�飶��b$.C���4@���_�;;!�Ue�/�1']����>M�������J�fHE?��F+����Y�V�R�I={q�3��Ța�rG�w����̆�E�eyF���s��[�9��&��u���hXݝՂ����_x-dn�>��V��5�/r�CKu����S6��U��#�C#���?D�sW�)�F ��̛3�=S�}g�Ap�Mַ��a�Z;��Z��)z&B���9����U9�/ot�����ܽ���!�	�k�O g�V&ʒ·�{*������;2�:HԫC�,��r�Y��@����0ں]Ǯdc��2�I�=�����Yhv7�'Ilz��d4\���H���畞�v����2���K�eBD��Vú:�FQ(K�V4���[��G#e�O����@�MKw�\��,�<�8wz���`(f2F�f25=���a��q�&��'�	s��C�F�X�N�cI�?)f��5;>Kf�����g�!���:ˌxè�k~�k{O�kbI)4��>4���ҋפ��1�H����,���x2$����zǏ�X�u$E�`�����$�zz��:GӬH�H]�4��b2����6�y��k�h�4y� ���-;�GqT�G�&���w�C�|�ޓ��dk7��&;r���c|U YMb�{u&4��p7P�_X5���Q��{�s�$���$4w#���V��axN�C��ݻsu�����`�P�"��1a�0�';�ap2�W���0V��R)�^��Ç%7H�̃�@�K_�R�>#�άnU|�0Ѷ��}�|�!d���+c�W����9��2h�Z�#��b��Ftbo�@Y��*��j���������8P��R�S7���3��Q���G?��z�ɥ㢐H�^�Ž0ٝz�:=R!����^fD�\�ҢH�#�O�[<��HM�$K+�NӠ�~��X"2M�D��	ma��;R�(s��G�y��4��2|��#�r���$õ$�J5mx��0���$*�a��:���S���S��H���"��W��EHvP�O�~H�֊�p�'�-m�����X��
Y��V�'ł�8+3�;�;/�oR�u���h�;�,C�aKN�-����@���yӥv
�K�q����� -�!�ֽ:�P�
̺r��>�{0���r&4FW	��^��.���?�߸�/�IT�뫾�c#�pZ���^x<����̩ʭ���<����{?+�� ���T���x�d� 4�rY�3ʏS�*�o�
��;E�VY66����Љ��c^��2�����<�k	X֒��M�O�P����ճ�s뭨i����`�e�=ޣ�����qѺSr>\�I���tzl��r��~�<
��{bg�eY]avN1�0��$C>���۳�Ogmi_���0:'��$�E�>Pԡ�����:gꡎ.��~�~*���*�%�G������J�'rS�I�;�y�ɥ&��$�@�R�tF��<`�HDӾ:z����ɚ�L������H���5��)C��#��W�>��F����<V�����r*�u�v4�o�P���E�ݘxi��m[ �Lc����5�{B��nNs��O䪷��M��L`�� ���,�6�}\P�=�Z#��������ɻ�gZ?f2�~�ΔH~�o�S!sv�fNߥ�|��}����|�U�'L� z�n)~��3y�r��d�5,�n����\h�Ԙ��(��}��Byҭ n��hEk���J)��?T0�� �(�7��o�]�2ݱhec�EbiF���!Y�G�����2��8 b�\w��!�vy2a����|nPϻ�����F/��~����:�u�ݡE��a��kJ�����E2�ZP��E��l������D�7����@�e��cd��m��_�mp�F���������
�mQ��v�fQ��~V����/B��d��&�j^�(M�k3��H��IY��ښ�`�+��u�C��V�C�	yy'�'�*R��ܼ�N���2��@(b�كe�DEx�9ў���E��O�a·�'�{������ZG:S2���%Wqp�P���N�R� ���{�	�V"WR�o^mC��\�^����cD4;�[�XѴ�]�NT�=)��(;�Uw��Gh��P��|,m��Ԧ _2��	9665�s��SK��u'x�|{c5��˪�I`�φx�\�zC���]��]�R��t��P0<�[Y�	�J2��Z��˵f���#�%B~P�֤~����o���xQߙ4�/P0o�����y0���c)��}E��t�"���n�A���B�X"���:h%����!�Q��0��Sh�'�hv����l�00�Uv���!>����'�&��=��ox�����M��\�{RAJ�Mt� �%x�l�6�?u��ݬH�;a���HQ��~36�B�c�SG�8�TW+xP!%}�v��/���[LZT�>��ӓ�d�'��w��VJ�ZD��ıW�ax`~	n�))U��/\+�pJ������m�a\~h#X�Y�Rǁ�#h5tZ���|6®nZ?�4�\1D�� �>1�M2Ђ0�o�HS}���r��>�M$=2��%�*m��OXP�/J�'zBڢ�QL�F�u�����	����r�C�v�aO�]��J?�F?�(_[,k~�"�}=�d�ȥm�Q��uH7Ep=C��3��غ5g= �1��A轝��GxZqR��$�e�f_{WW�6��Ze�n�!��8`�dx4���Ht Lϑ�J�K��=�B;�[�쵲�7Kk~ؚoÕ��c�h��Ex��6�5��>\�~Q�����\�$����jPSs� Qyo6w�����7��v� -�]��,�&~}9���®�_�cc�5�pc|F���|C�1i~Gu��������8�:��/�_t��[��U���ʧ k�+j�V�ž�%!ˎ�)"�]U�"��Fx!IC�Yv�������b�p�O�gGn���HMX^�l��uJc0�a�ҽV_o�K�_5I�qz@�i4����eAE�̣���>��j�?��o�R��E�P��;'���s�n�
��Z�Ih�oUtUG?.�v+�Q��H�����K�0��i5�fR���b�#��n0H`=<�H.)" D��W�)ɳ�=J���w,�J"YӰ�S����'�OvnY���lz#�u�ܛ!5�C��*Q	�K�rG�#D[��� ؜�@q��e��p��/�ոշ!L�f`X&����&Gj�%�;�|>!�=vR��������uH�i\7<�SG�^�;�Ӽڋ[�	+W*��O���
��^?V��YhS]<��m1��\�`���B3iQ��6��p����m��){��Q�$p�U!��i��U����:��h��}��w��)�&�a}�|U]����CqXΔ�3q ���7�>��j,�����[����c_iu)'�h�Q�L��@�(ߝ��������q�� I�Q�a�kz�35"��@L��X��Q��o�˽�y���I%�j�$��4��ؤ�\�`͕�jf3[���@�j�I���	��\w �.�ԏL|��]�@j��Eam���i�Q���*���@�LS�Wf�+ ���QÂ(�|�^�
�GW�*q���t�ǤS���y62��^ο16dA�T�$8��ˊ�e��� (�W��rm;�q��s��ɶ�1�o��"��=T�I4tN�5#��x����V��q�>�X9�[�� �D�z� q�~�k(� �qYGo��^�!���d	*v��C�u.���m?A��P���x��4�sje��m~��񖝮��_��O��HОɓ�׮�YZ�0Fk;$��8���iB6D�}V[��%��I*�CO�6r��4i�
����_E�N['�
|AB0P�+ٍ�|���Jinܘ��9�G��4�S���(O�������6�=}���E���tPK�,%�g=��\�O?%�>�|���P),��h/B|�PaK��
/�:J���N����寲1Z�F3���'����u1zH#�&������8襯�G����vJ��92A�f��$�Di]��43���i�j	Z]�yT�lp���sYiȰ���� ��)UL�}�ݣ��ꎳ�'����¹E����W�0���>�"�z/=j M切���dC��~�nr߀�^�s5W`�sv��"eHl�KE��+1m�S�{-�S�r5C���^(5�-7�	g	|�R�N��v���v�����^3�b�6chD��7%h��ݙ���UA�׋��/�\W��mhv�i�W�C�'�c�F�h�A�u�I��wP�pb2\,����Ή1���Ŭ����[���1&�r[��5�x�m�	�v᭛��pN�/�<��?��é�
�"����æn}����2C�Uy�c�ʣ������ւJ�����8Ssm��5��YD��*�^����z�t8�������M��	���y���P.l�/��*}��N�ss�M %�i������߰!�/�y�[�ɥ��D2���z���ޱ��BQ������DT=��X�W�(IQB��&���ͯ!�;��v����47�3��(��㑘�LXw��˜�>K"��s�l�����\��Һs[���5���k�v^�S*����u��)(BG�ʘz�>T��ln��G�́T�I<�8*���|�8�-vE���j����/�6(���R!T�>�+�}A4(kK�.6E��0��<��wH2 Ms=�IqDEO�?���i�t��˂��#����l���
x�;��}N�*��"���0�~~���Q��=���F;�"��������/����j<�T٤���b��K{	Nx?��]w�5��ʭ�q���1��FFӳ�r��Q��ܿC}�*4�uFZCf|�6)��\^��F<�r��*�����'����'W�� #1ٺ���o�*[Zyk�#o��*r�M��J��1hh��E�m�7�7|W��ȼd�25��F-LǪ��Mݏ���Q� ���i9��O��x<��ִ>�#JDZ�a����#\J����IWD����N���6��}-4u:uJ���٣�����	��KA��]�=�(�^zE�v��.^�q����2���Vq�����(] 6��9�����4�K�>aU�e@Hq��e@0/BB��T�'%�.�RhjdN`�:4ڏ �����V���`$����za@�J�>N�w�w��껡l�VoeJ�P���N���m���#K�{�%��G.:7rK�n�p �gX�G���7ϋ��,���M)�e9lnΔRZ�A�H�gyn�N�*�<v�������e���:�L�u��c 5�DD����DtE"o��I���"=�d�P]�O#�d���g��[y"<Ї˳&hT+!�ȗ��Ե0p�lF��(D��s�4^8�Xj�'rV�A��CG-~F+bn��+N�B���7l�
QX�6 �-�H*����M��\�g��H�nU:`�7�u2���j�|�s|��B8��nEx
�Ve�K��O)�"�m��W��|�G<
���'�?Ía9hdON��d/a&2��4ҷ	�/�,��N\�mM��a�*y�%��_`@����O�%�29�z�2��ν���Q�1*�S���|���ø�S���S�y>sp���h8�:xSm��Ʌ�@�璺%q4�ȁJ1Y�"���?]����=1�V.����k���<b����c���e�*��D0�����\B���+�;�Á^l��Sd���U��;b��!F��%mR\����kɞ���ꖪ�	#�,��v�E�Kzdi<���<�
zmUqm�ʅG?�oeW�$���Q�D���G\�j�?�SҙXׂc�U@D��O���%4V�I���m��#!�PτUIr��F۸	�a&h��4��T�x�:)~`�WH#b�tT�V�p31]�r�]��h����<B���Ě�)1���=v�	�[N�-�9���0nH���_r�H�莌���Ii��d;F����[���\(p���M��`>$L��Ú���n��~�I��6�� �%��Q�GY!�H�_���s�Z/c{ �c���Au��y�`O��?��2]���O�Z�iu���d�OY�P�RZ�Fǽ�E��F���TXBʀ�9/#Ԋ EѸ��u{��7	���w��ab N�T:	�������w��ǈ4oN����Hш���J߄����錆Bnmߺ:�-�̜�q�F�� �	dή�a��{�2��*}![z���6�I�H<���eE�}ߘ �mD׋�Q��B@�2������u�p��F�[�M�[�A��q8̤�Ҭ�t��?�'7�.�����Um��QA����`t�,��o}�o!S��T��6g�s��/����M]r8ާ+�{=n�;����`��,�����u1��3�/G�>