��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�����g��y�(.��H�^���z=ͦj�P@���I��_]�E�����U��@�iKAUu��z��}Kk�4�m�dC_�0w+�͹.a(:��D����ɿvw��s��=��PS?�8�\р��9ꌭ���:`��E=��8u3 ��;��\������k�@s���|������)���J �ꨣ�҇�6Q�?����G�����d�@hc͌o_� U���"U�4��ͯ�>���l?f�7h��z�U�]�\in�+4��l
[�W�*�鉪G��Nj�lzR�5�bV�����2���+�+�[��Q_#(�0h�9V�C��N���P����r��-���s�vw+�j����_	N���h��TY�j�N��x�8fy��_�OFZe3�e��CFY���@���$-9��wD��I�+�=�K���mI�>��D��>{NK�cM��e�Q����Tֵ�����H�)�|B��t��oXL��@��3�;F%�i���6�=���pKn�_�9^��3�fz[��_a���79��@b��n���,��{�M��EL��蒠�7Dr}u�bA�3m����{��Ȫ���4l�A��?v��(2N$���Sj[�=mm�?o��И#kg��2�~��Ui���X���dM⎷���4���`��`j`�A��xalC}C�?�Ło}�	ȭ�몽y��)x�ɏ��yx���9p]�\��DL+Xޙ��T_�d�=�C���)*9�A=;I"&d2`�Ȗ���8��t�F�.�ӆZe7�~*B!շX�UTc��O�!�熕j�h_��*L�K/�Һ���1��W���ٖx��ꐪV=LZ��(ҭG๑Z��e!x)�{>�n}��Ԓ�Z"0:������z7;�,I_K�Jl<��pkѨ�4k@@5Q�r�<�p�ZD
<Jc��=�*���.nH�,�!ws�ڲ�[�L��}�({r�+���y�|��P&���4B�VK�-�SE�A��K#��(P2l$!(��h����Ԥ�_�y08��h���y�e���H��Ũ�4����H@�떞_��d4�AY���zHB�fȋ�!�m�:�P�b���o
ȫ'q^E�	2tG���\ǡhi������ּ�!����!:]
.<1}2���6؀�	Xd����&D{��c�1E�RDY�W[ قs�c.)��M�ε��?;�pI�/�bە+}&��<Q�/MP}����ܥ�
)���M�{�s���j�A��-�c��ȸ���V�J`�f6cm��אD-�MՆ�[cL��/F�V/�b|�@���<pt\�F���,�f�Z}�~ߑ�.	����q������M��u]�@�"z᳢�m�ͥ�ҵ�YP4eY��z;��d���O85�4��+ne�H#�z���$���y8 Cu^�Ĵe�H�O,��"��V�Gٮ~F8��1S���h�����A(9x{Ӯ��� �=�?!���o~��8����2�/��X�y���+j��R/"�@\)M2���ɓ�t	;ɣ�]o��o�`��k��
@�~�	�P<N�e8��&t�t���� ��Լq	���RзޙE2׃�pP�a�?_L>�qڎ�CYu^1R��*�?�!��"5P��$hw����}�ܳZ�Ȧ�=�Sw��(4�����)0�©i:/���L����Ms��_��\"���lݽ�s�k��(�ES�u�
{��� �{��
�u�rx�;���,AlӀ�^�&P�G�S%>ba�.;0��WR\:�~��o��  <�-�V���
프 Y�&m��<Hy�	%�@9J��/��70�i�)o��U�}�}�17���Ql�|���E&ҬԨ4!�O�jm�,0��&��$5"d�\fEd�P��(wd�Lח6pUc���6�T�QM%�%C>�=����q>֛���L1!(��X���?n6{jc�z�"Uc�`\�=eG�T��W�����S�
I�]7��qei~z�����E�5�2*�"m�
�vT{�MM��E��V��A�hz�zU���U]nRB��RD����������L^Pi�����:��΍���wC
�iP˦�U;v�S5&� ��OA����`�z���ȷzJh���"��o�`�Β���^|n���,�Vy���.��_�1�?nC�N���ߛ ��fpNW�La9-�jBp|��H���B%T���ѽ�d���2�MRW��ꇗ�Ok	�AP���Vowx\�Reʅ�4�$пn�K��A9ҏ�5���$v�x�t����>��!�%�N�g��Ϳ�;�~�Ș|؏�5�Fg/��g���������l!f�ؾ���-���ۈ���XB�:�{o]/��d�6�q	c=~������go@����V��-����TCo6p�Jz��*J���Sj��nbZڛ���s{n�~A GX�%?wbe���r{GȬ���C/\%S}0g�@��½7"�O���XV��MI���%�6@��$
� ��|� ��4��mB�'�D�A��,�E�73<�|��+THh��Ę�vU�����^Uk������N�<K6$ߙ;��Q���Y������#�[7�І2Ǚ4�Vh��B����N��;H֘#��r��M͑��8r��P?�D�0��N�&TޞуQp�"g�P&��÷���2}�F�+L&��E��5��77Ӹ�y�<bh²i&��;A��Ӂ��q��?�'�q�S���<"�X�)0�hK�#���e���k8�g��n��nLG�Jn�nk�"�����^�Ir��q�H<|e�\�<�@�f���ґٗ&NmN[ji�XhY��������͇(<��<p�1m/�)2)��Qcm:��i���Ƣb�f�c��$1ool�QzVN6!(��J��vM6S�����H���$�
�S)&�he���ه�A��%���������;��10|�P{��$�x�sG��&�n����=�eU�&I�.�j���X~EF����1�/ʭ{��2�;�I�r��Iw)��K;�����ǻ��R��-�>�T�!�?�U M��1"ō��ife�[������Z2'z�ך.y��d2�Q:c���_'Z�'�3����[�������
���.��N�n���D%n�E�/���WI�g��� :��C�F)��Ҵ��p�7l��UU#Z{�n�ow� i��88�D+�kc����͒�Q��%���b�E��E���o������S���4��֤q�&!�<�����Sɇ�|��-Â��� Z%���%�:-��t���HV�� �}P�Mq{M��lo�ں�!��v?qR��]��f*=���|���]&w����*\�.��7d�S��}yϑ`�Z��6��X����+�g����l��s���ⱦR����Ȣ$��q�mT\ˎ�z2Z6�&0+�M;��S����}�
ށ��x!���Af��v��V2ݵ	�]�i>����m�~_����ژ�N�IJ2A��/>i��F�� uf-%f�V�����Tq���	�͆j����x���,��]}���@秐�o��$Y����<��oTx�����p�#j����m��ys3��?����n��K=3�HW�D�)5xE2�ZMyԗז�2���?�ތ��)̤j�5r����m��k\�V�"'�鷥s��U���q좾uʜ�?��Я�Q4����-	���[������q\G ��Mx�,���D���1�Q�'�����i��D뼮є����}9f�anuP�S���J�m@#�m�2��5�����t��\
bƥ�b�֌��Tiү��{����y8����Y���H��B��6� '��8�c��������� ��wO�q.�S���o��QACR�&�e��q�-��9슨A���l�Km�&�����q|,���܆���(���Ң��9�&F�F�.�aRi^���]�9���zI�ޱ�K;_$�ƭ�@U��Ѭ�»�A�$f5��3Pc�d�����H�c�,]�6+C��1w�Au�k���O�CS�����H<Gz&�.�v��g���4ʀ+���O�	��+�J���ե��B7��.[���5�<�:q���,̖j��"p��J�E
Fג�����������%��&[{jcȆb��ZH��Q������I��A?y�/�U1v-SF+���	/�㱫��p,�I�t�������F�����WSR����IG-Nģ1|�E�$M8Ƌ�/G�M�|�	��{���L��>�ǩ���O�X^����h>W4�Ĝ��ǎ�����R�oh^�f�k�39PxL��^N�A�5��zL� �s���+���@Y���M'ڊ�(a�;��.�ܔ�Mۭ0׽X�V��z��d?��~:݈ƔxA)Hq�<��5HC)�R$�m<+w�c&;���#`��",��&�w<}2���sE�
*�!�Ă��T8j咏�i�_�(�+d�߸ֈ't�1�N��Z_z���"-��_���y 4ѓ���H�$Z�!J��L �J�"C����<���e��y�-�R���Qb�v.p����!��k�D2�PB�܈/{+�L�u�88T�l�מ�c�X7ߴw*��5���y�`/��3���Ėf�Q���z@4<3cRujW�%(�)�����l�O|U���f���5b�=~����x*����u�cZ}�}B<���iVTd56���\U=�}�9���d���jt�ɢukҤ��	㝫��&�c6��[�l�/�L��ĳ�	.;JT�@��$��u����� K�8��\����V�J���8�������.����n
��o<�Jeu�v�*��7�ZA1�]IGP��@��$mk��cV��	� ��VDDi.Z�,U2x�c�c�5�\�q��T��9��Xz��oD��D�&�����EԥM���qb��Ǌ�Kږ"2���4�l��|�:{m��̫?��%Ҽq�����g��r���@�]��A���K7�8B��c��؅�l��݋����!~��o7�ι�wQ�EP��^��D��=}�y�9m%��*�.�]���_�}�m>q8������Ϲի����I�e�ܹ�uh(ށ�I*nQ����ntXT�ȟ�Yp�H��EH�!�:�goD �W_H�z|�V����f�C���r��CH���.Q����Lr*y�:$鬕���Q��{w��R�g�#���,�"���� �T�v�V�3��j�]2�@�X~5|g1y!6�*�E�ɦ�x�٣h0znOp40@�_��y����e#â޿���,��~� |��6T�l�<f�V{�sk��L�Y:�/U�J;�%!c�-�	���Z1دN�^��1�x=�nĖ��N��X[����jO옾R"ێS���V(�$��!���(=&@���w�'��YbUfvz�$��\)`"6�:I(_؜#����W`��%�~d��j��1�u�&P��%"����%u���qs����ll��$�^�ԡ�d�S�+���?A��#xz�8z"%��4Y�m6$�E�p�|��k�;9s��u	TW.�QS��d�c�>��(��Z�.I�@j-��+�*&)r$���g�ܶ��r�>,�7�D��!�����V�Ԇ�W��a��5=���X����T%�S��������!M&��|�m#c�LF��΂�K�,����E�8b�D��d6o$��ߗHc*��ğ��~�5�J�8��x�^��-�b�!��,�</�g��v���?��\���\���קo�4')u���v"Fy���+��G���΄��5R!d�/G�6��.o�7�:N�"�%�r��UsHW�N�*������e�c�x��N&aZ3�2F��\�����N��OoJ	�ڊ'��\F�4~T.j�Z�tV�xʉ}��e�1di��qU`hf��[�L�ߡ��@P:�6�Q*�"h�}5e��	��`_,Ǹ���ݚkɖ0��&�i�7����bq�;6�, ����� _��zMq���.�F���-����%A��'�����K)X@�:�9���
�豁^١/J��Cf�2�+DC*������ło

X?�f=���mM=T�:�Z/���m��9U����.��S ����u����P
7��T�u����2��F^4t'%T�5���[<����w^2�>.M�5/�iA��!'��kY;�{����0�)	���+@)�"dkl�*w�Z�W2��Xw�z�N5�(�����0S�� ֣�(xOY���ΩϢ|��A�e)/�2��A}�k��`�~c�
C�B%~�(����K�������O�ۨ�k�e*s�\>��d]��/ٵ��P�%X�d�ʗ����Ԟ{T�2��B7���w��>��������9���@cP�h���6*L�-k�*~�F2J�f��XS�)w���4�8�,'��P�6`35��y>%K{�olMf�>����9|ˬA���1��������������T�z����0󘈞ʝ��LkΫeB�p�r���u0!�B�y�E�
I k�F�j���].�d/�c�w�ْ�S.���E�O�YY�����z�%ʝ�8����QկJb2��|y/+k XT��}E|���~z��?�Z�� TVvek*Ub s�"�o
���`֐�np