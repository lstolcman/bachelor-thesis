��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�Ji��R�*�u{"�sdTE|���wkSm��?L<��G�»�X����B�f�H���͊�6NB4�)ư�X�K�'��T�0�A�%٤ޮ�Ѝ	��yH���{x;5�
iݤ5��2��)|:>��ǎP njL����a�#������x����У$�֑��v�ߢ� �zWd5^aR�h��foF�9y�jo��;n(�
嬆:���5q�v7����a9ڝ:_�
)3�!�\cN���@U�z�*�f�p��G��4EX����L��̣�Wh�tKE�TKW�g���%�+N�B�<�~�q��T:88"g���K���#%��5*�:�P���.�l�T�w��G;C�{�����7�;��F![_��HU̥m,�A���^��#�������\}=���z�4KXh�|��)�`�9�n�E�s��:���W�ti;65� �#�sJ=Kf ]KF�J�1�Nʼ�\�����W��;���E��jG�]sd�U�4��z��^�>�,��}a��*�n�I.�������}�Æ�O� �֙��#���Weܱk�F6��DRL�Ǧ|DQ����[��au�ƿ*�%�ƈ�^7w�6�������Pkw���3��Ά�q��Ca"�A��G"���Y�v?
��$���4 ��x�?�0
x��]1�I͸-\��!�Ц��w��7��6ކ�b��G0�nG�̝Q ���?N�E���b��i���_=Bu��?��19��89j([�������yb��}!:.��Lb��O�u�%�ع�u�y������3�5k�����A�Y�j���&h�9`�/!�ޛ��f�&&�z���;ca�G��]��'��t�H:��a��8{6����~��)r�`��	�>�? �'���2ڦ���13��<��NK�seG.+5�m���R̌��&���t�$`��F�]T�0	ʬ�1Y�*Z�٣%����]�z�oWKk�0� *�OI��>�k��y�uʩlޕE�p��#q&�r%��hX�Cy���Q�#	6�2��OR�"�$�-D!�$����yR}ե�Z+��3Y�X�Zq�q�_�Fx�B��o}v���4=��W�<�嫐GET(WXt&�Tҳ6�m�VE8�uL��@��^���d��DA��oB����F�ЈӦL�)�k�� ;��߱�q�k��go�UL�w�V���y`1~�J'�m[[���[09<��Jo��c\˵s��	�VC��of�0�8m�m�:�MѴ�c�wY�3H�KiDB*/���N�+�ľ��_��A���q�}�_q��a�TȃΧ���w��2x��i=p� ��}�?�z������@�̉>��4��p�^��"ri%#�7�v�/Ĕ��80J���
8�1���
�f�8'��������b���,��i���08��;�p����<R��f� \1;i]�e��~�h������3D�Ls�z&�*_�����Ho̚J�f�"3V�V'Q��P;$�b�P "�M�oc�q8ܬ_Dykvg���8[���hC��I��oS\w��|Mj��������S٩�4�i�����+����l��碊`t���m�������|��L
Ы([v��듧$�����/�I��}>�k��l5�9�CK���c#��#�X��TŌ7�����p��ek�I�����P���W���l-�͑&�X`(ul
���4{d�K���ޕ$�U�Atgf|�8����h�2p���d�l�^�Bhs�Q'�"��A����sq�A�"� �S^BGgs�%�a��P��F�7s+IO��Q��Y��,�ZwڑB�� Ξ�
�}k�3�]ٳ�lL�U�d� ��-�R�@�H�C��� <ѐS������7�	�뻤) �!��y��� �s�i������͒��d�S��ΠG!������P�6慕4�R�w�����|LA��'w=A����T��.	��&�@0��2�;���ܥ>��� <�i��Fv�i�p��V�&(���T��5�Wr5fb#L<����a�#5d57�����8iX��B�F2ʸ�%=��H��~	�}���6���A�sًV��ƉM݊���䝨:B�[�@2dU�`P���_�� ��1$$���	$��O�t�1�Uk�.�;<���
�!��8�|��.U?��0����8��3�e������~���Z�=�waC+��r�����2%�M��<��T���y��Ae�f� ���]`k�c��l�$堤/�k���8,|��i�)o�.n�8�������/X��a9�7�1����������~���`^��a��n�ʱ����=�=6P\��M�V���f�)�0ۺ'bE�/~���h�MݲH
X6����*��ҕoP`�H�Ŭ�B`;��eH����Pc��b�W�h�����r�&˦���wչe�P���GϿ7X��[�!�6�x�y��=�C�G#��S�E�g�J�pm�C���uR�0�Ҟ�4�t[{9(6�*�IkH
��Jf��L�֩��狋?��ܟDǥ�;�w��	�S��/Ȳ��j)*�hSL���);��/Yp����˶%�.���%T�0�:V�
���	��7���	H�����(��B;$����g��2
���ϲ����.;t�Q����>�bY�3rB��o��ӄ�?�c�>tg����f�EN���޳��9�A�e�ɡw\t�kP�P㡶��);�Z��X($��CUL�<�;}�$�.���	�;RƷ��y�=�^[S@��N��^+P������q��L�^�6cYO"$�C��>�‮����m9��	�� Q����ŕ
�!y�m0��g�b����%ҺI�t�&e�]\��Fw�M'g��!�H�69W1��iO���:����t�����Q��'M͢P��h]�|�����v%Z��C�\�#d۟����7r<�=[���C[�4M+��Xo'7>$�6� T�0���Ґ������h�T��#�Շ�G����F��H���s�,q����7�?ڻGJt�}6��R]�^��,%�~����d��++zӄ���Y}n�#�����7⯄��`=�s���PS\���S㋽&Ȫ�H����޸��W%:�d�Ҹ �΄8�J�ٜΟs�M*�!k~a �tdĜv�*�z���3���ݷ�Շ.�2]�x-��ȕ��ן�d.�O8�z�{���u�t�T���U=��L���2�*�/,4�����e��Q9�&�ә�E���F 5��ķ[`�t���TL#��G��mQD�ܱ �������n|{.�,�ֺDo�N��
ҧ�����{J9�Yz������y�x��7����Lg�٪M��yThE9r"���$ΐhp�6���;��}$����'c��)�K��J*��
��Q6�ۋF�|�GcH�s|S�Qξ�xG|rQ�է���4A�9���F2�rj�vk#ْؓ1z�Pr���5]6'�*i�A���NS�6����< R��T�n�\�w[��|�/����&�F>x6�7pn�*.+r ʎ�݋ˬ�Fl�N,�'h�e�8������"G�/'&�x�ѕy>(�em|f�k1|���E/xvV�a՘,����d��}s疢K��>5�{��(�'O��[���`]F��F>���FRJ����逨Bsy?;M5
����Q��.�*�3��Q�Bv:�I�K�%4L��s��%g�,��E}?Ԏzk1�TJu�Cc�M�~H�W�:=�4��P�9"
�˔�MfUSFl�������%�U�C�Hƛ6�8j�.�����S����؏l>z��qM��|�S�h�XGA�����/#	I�4nS���m��mH���rj��.vL�AfC��EYYa��|*�Vy��R�2y6��S1�k��/�� ������g��t&��_�xs��\��� t�_̚q�8=P}����+3��!��&� ƖJ�������U�m�<E��@zU��}ᨀ���ä�ҏ&��n�ݛ��L��(V����
	����a��pj�'�Ӧ>BԞsz��[���d8Vf�UO}Ϲ��St����಄��cdXY�� :��^e� ��jw�G��M/����N���3���kh6lސ�`�M��o��$COC�0�A�=@c�c�f��[��9pV��s���|�Od�[0ͫ��s�j^H˵����Psa�w�N�??WdF�A����