// megafunction wizard: %FIR II v15.1%
// GENERATION: XML
// fir_second.v

// Generated using ACDS version 15.1 185

`timescale 1 ps / 1 ps
module fir_second (
		input  wire        clk,              //                     clk.clk
		input  wire        reset_n,          //                     rst.reset_n
		input  wire [25:0] ast_sink_data,    //   avalon_streaming_sink.data
		input  wire        ast_sink_valid,   //                        .valid
		input  wire [1:0]  ast_sink_error,   //                        .error
		output wire [31:0] ast_source_data,  // avalon_streaming_source.data
		output wire        ast_source_valid, //                        .valid
		output wire [1:0]  ast_source_error  //                        .error
	);

	fir_second_0002 fir_second_inst (
		.clk              (clk),              //                     clk.clk
		.reset_n          (reset_n),          //                     rst.reset_n
		.ast_sink_data    (ast_sink_data),    //   avalon_streaming_sink.data
		.ast_sink_valid   (ast_sink_valid),   //                        .valid
		.ast_sink_error   (ast_sink_error),   //                        .error
		.ast_source_data  (ast_source_data),  // avalon_streaming_source.data
		.ast_source_valid (ast_source_valid), //                        .valid
		.ast_source_error (ast_source_error)  //                        .error
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2016 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_fir_compiler_ii" version="15.1" >
// Retrieval info: 	<generic name="filterType" value="single" />
// Retrieval info: 	<generic name="interpFactor" value="1" />
// Retrieval info: 	<generic name="decimFactor" value="1" />
// Retrieval info: 	<generic name="symmetryMode" value="nsym" />
// Retrieval info: 	<generic name="L_bandsFilter" value="1" />
// Retrieval info: 	<generic name="inputChannelNum" value="1" />
// Retrieval info: 	<generic name="clockRate" value="1.3" />
// Retrieval info: 	<generic name="clockSlack" value="0" />
// Retrieval info: 	<generic name="inputRate" value="1.3" />
// Retrieval info: 	<generic name="coeffReload" value="false" />
// Retrieval info: 	<generic name="baseAddress" value="0" />
// Retrieval info: 	<generic name="readWriteMode" value="read_write" />
// Retrieval info: 	<generic name="backPressure" value="false" />
// Retrieval info: 	<generic name="deviceFamily" value="Cyclone IV E" />
// Retrieval info: 	<generic name="speedGrade" value="fast" />
// Retrieval info: 	<generic name="delayRAMBlockThreshold" value="20" />
// Retrieval info: 	<generic name="dualMemDistRAMThreshold" value="1280" />
// Retrieval info: 	<generic name="mRAMThreshold" value="1000000" />
// Retrieval info: 	<generic name="hardMultiplierThreshold" value="-1" />
// Retrieval info: 	<generic name="reconfigurable" value="false" />
// Retrieval info: 	<generic name="num_modes" value="2" />
// Retrieval info: 	<generic name="reconfigurable_list" value="0" />
// Retrieval info: 	<generic name="MODE_STRING" value="None Set" />
// Retrieval info: 	<generic name="channelModes" value="0,1,2,3" />
// Retrieval info: 	<generic name="inputType" value="int" />
// Retrieval info: 	<generic name="inputBitWidth" value="26" />
// Retrieval info: 	<generic name="inputFracBitWidth" value="0" />
// Retrieval info: 	<generic name="coeffSetRealValue" value="1.89907364531E-4,2.67905072965E-4,3.06622826868E-4,3.02119101944E-4,2.56217153567E-4,1.76173836546E-4,7.36781004787E-5,-3.67179960185E-5,-1.39562137948E-4,-2.20623519929E-4,-2.68897320107E-4,-2.78205763036E-4,-2.48140073812E-4,-1.84162038471E-4,-9.67981167877E-5,-5.12337876497E-20,9.11080208379E-5,1.62748844873E-4,2.04855412159E-4,2.12843665209E-4,1.88434049417E-4,1.39308037539E-4,7.75913677805E-5,1.73843240496E-5,-2.82313758038E-5,-5.01339910233E-5,-4.54313927947E-5,-1.85152538923E-5,1.94474703511E-5,5.2642663598E-5,6.40776434848E-5,3.97928044135E-5,-2.70143525424E-5,-1.32873538917E-4,-2.62765964366E-4,-3.91247750828E-4,-4.86108142638E-4,-5.141901471E-4,-4.48500105783E-4,-2.75339595489E-4,1.05514097046E-18,3.50369131836E-4,7.27752329471E-4,0.00106855008446,0.00130280847846,0.00136624533675,0.00121322353325,8.28381102836E-4,2.34558587079E-4,-5.04975270314E-4,-0.0012912228806,-0.00200120881138,-0.00250565372767,-0.00269023840495,-0.0024771949253,-0.00184350362909,-8.3212085516E-4,4.4654659123E-4,0.00182433977331,0.00309587922358,0.00404770259427,0.004492078925,0.0043003649969,0.00343031598861,0.00194220984205,-5.11278586565E-18,-0.00214417217498,-0.00418118467761,-0.00578827239929,-0.00667859638691,-0.00664961136729,-0.00562235533085,-0.00366459502997,-9.92788865912E-4,0.00204916572168,0.00503286810374,0.00750491718131,0.00905484302697,0.0093813997159,0.00834670021565,0.00600887256799,0.00262667940388,-0.00136647369647,-0.00541707308275,-0.00892790710392,-0.0113458605228,-0.0122482090293,-0.0114140250417,-0.00886887302752,-0.00489447371296,7.91665901847E-18,0.00514257609598,0.0097910024104,0.0132403691225,0.0149301546908,0.0145343932386,0.0120205317221,0.00766672143646,0.00203321556298,-0.00410962789473,-0.0098875334685,-0.0144479407165,-0.0170868570053,-0.0173578944498,-0.0151465249619,-0.0106973119078,-0.00458861109969,0.00234299658056,0.00911863528157,0.0147571775275,0.0184191102281,0.0195328678732,0.0178844204258,0.0136559985834,0.0074071724391,0.0,-0.00752164038269,-0.0140814014084,-0.0187268178057,-0.0207696139655,-0.0198890102481,-0.0161823273961,-0.0101548608373,-0.00264995070515,0.00527093008993,0.0124807506097,0.0179498831329,0.0208955190185,0.0208955190185,0.0179498831329,0.0124807506097,0.00527093008993,-0.00264995070515,-0.0101548608373,-0.0161823273961,-0.0198890102481,-0.0207696139655,-0.0187268178057,-0.0140814014084,-0.00752164038269,0.0,0.0074071724391,0.0136559985834,0.0178844204258,0.0195328678732,0.0184191102281,0.0147571775275,0.00911863528157,0.00234299658056,-0.00458861109969,-0.0106973119078,-0.0151465249619,-0.0173578944498,-0.0170868570053,-0.0144479407165,-0.0098875334685,-0.00410962789473,0.00203321556298,0.00766672143646,0.0120205317221,0.0145343932386,0.0149301546908,0.0132403691225,0.0097910024104,0.00514257609598,7.91665901847E-18,-0.00489447371296,-0.00886887302752,-0.0114140250417,-0.0122482090293,-0.0113458605228,-0.00892790710392,-0.00541707308275,-0.00136647369647,0.00262667940388,0.00600887256799,0.00834670021565,0.0093813997159,0.00905484302697,0.00750491718131,0.00503286810374,0.00204916572168,-9.92788865912E-4,-0.00366459502997,-0.00562235533085,-0.00664961136729,-0.00667859638691,-0.00578827239929,-0.00418118467761,-0.00214417217498,-5.11278586565E-18,0.00194220984205,0.00343031598861,0.0043003649969,0.004492078925,0.00404770259427,0.00309587922358,0.00182433977331,4.4654659123E-4,-8.3212085516E-4,-0.00184350362909,-0.0024771949253,-0.00269023840495,-0.00250565372767,-0.00200120881138,-0.0012912228806,-5.04975270314E-4,2.34558587079E-4,8.28381102836E-4,0.00121322353325,0.00136624533675,0.00130280847846,0.00106855008446,7.27752329471E-4,3.50369131836E-4,1.05514097046E-18,-2.75339595489E-4,-4.48500105783E-4,-5.141901471E-4,-4.86108142638E-4,-3.91247750828E-4,-2.62765964366E-4,-1.32873538917E-4,-2.70143525424E-5,3.97928044135E-5,6.40776434848E-5,5.2642663598E-5,1.94474703511E-5,-1.85152538923E-5,-4.54313927947E-5,-5.01339910233E-5,-2.82313758038E-5,1.73843240496E-5,7.75913677805E-5,1.39308037539E-4,1.88434049417E-4,2.12843665209E-4,2.04855412159E-4,1.62748844873E-4,9.11080208379E-5,-5.12337876497E-20,-9.67981167877E-5,-1.84162038471E-4,-2.48140073812E-4,-2.78205763036E-4,-2.68897320107E-4,-2.20623519929E-4,-1.39562137948E-4,-3.67179960185E-5,7.36781004787E-5,1.76173836546E-4,2.56217153567E-4,3.02119101944E-4,3.06622826868E-4,2.67905072965E-4,1.89907364531E-4" />
// Retrieval info: 	<generic name="coeffScaling" value="auto" />
// Retrieval info: 	<generic name="coeffType" value="int" />
// Retrieval info: 	<generic name="coeffBitWidth" value="10" />
// Retrieval info: 	<generic name="coeffFracBitWidth" value="0" />
// Retrieval info: 	<generic name="outType" value="int" />
// Retrieval info: 	<generic name="outMSBRound" value="sat" />
// Retrieval info: 	<generic name="outMsbBitRem" value="2" />
// Retrieval info: 	<generic name="outLSBRound" value="round" />
// Retrieval info: 	<generic name="outLsbBitRem" value="10" />
// Retrieval info: 	<generic name="bankCount" value="1" />
// Retrieval info: 	<generic name="bankDisplay" value="0" />
// Retrieval info: </instance>
// IPFS_FILES : fir_second.vo
// RELATED_FILES: fir_second.v, dspba_library_package.vhd, dspba_library.vhd, auk_dspip_math_pkg_hpfir.vhd, auk_dspip_lib_pkg_hpfir.vhd, auk_dspip_avalon_streaming_controller_hpfir.vhd, auk_dspip_avalon_streaming_sink_hpfir.vhd, auk_dspip_avalon_streaming_source_hpfir.vhd, auk_dspip_roundsat_hpfir.vhd, altera_avalon_sc_fifo.v, fir_second_0002_rtl.vhd, fir_second_0002_ast.vhd, fir_second_0002.vhd
