��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�q����'��7�T�A&m��˴�:�u�����T5��Y�LN����]$j.Qw����F��&0�3�5�F�A�?���L�R��d��
�����8P����� NPZ8� 
�>��}Հ,Ӏ-6dvb8`�`I>;�g���:���H�f����u*��M�[��\��&���N��-Oh\k����x�SZ�)~�^�u(��=�W�%,�>x4I�m�ϙ����[0�l9�C)���$!��^�(0�����'b($	�rU�@/23�8�It�%)Pە@�z�Æ�������;>-e�dF��G�z,T��߷���1�@�	#��T@}r�z�v�{�{�,Z؝߉����r�,�G�����B�N#�_������n�[���nX<��9=�x��L&��F`wv�QU�.�f5�j�tH[��˚�1_aօ�33V�S�F�Vcu?��3?'�A�܁��Sۘ ƅ�Q��Fk����KMN�~�
;�a�6�W���^b��.�/O�\��8T|����ѧ%�3����_�%9-P���:��M�Z.r�X�֚�B �R9S�L\�ǭv�_�/#'�F��M�Đ�)ͯ���Ǖ{�����KE�u������;�P׮�3��ވ�l���������E
�Dc�����SD�'QC�~ݣ��
Cb�K�?���0��n��f�"c����9%���̭�k�ቴ�W��)�U�tg�}�T�|�5�<E?�/f+AJ�����?�Q�E�ŞD0�'7]Av6����2I��ͱ�t��r�ëvP|�@O/��;��[h��T5b"�~�&p���<�s���h*�WE�!��z`����� 1O �O��yy�u�sN�b�P�`�4�"Nd�rZ�mw���A����v+�p�r���<C�[n`�_V��U-�.�[5�S�[���$������lW�=�9� ��bF�ρ��Wlcc0"m>���ި�;=�E�H����2�Q5h�@�qK�̏v����� 'le�}�Gi
�'����N�#)�Ǖ �U��k�lG0GR�j,Ј�����<E�]޿H�L2��lpRv^��.��n�O-�Z�H��J�nN@=�R��j�PA�3���u6Iʖ�p	=^��X��4_
�[�(�ӹ��ɞjlb]����Y��M~�͸䛞���L�����9�:���D"�
�5\��@�C-,&��U���U�ݑ6?��7�����}������7%�j{\� ���E��)���5�7=�X����5mt`ӻ�4�9k
.!\�3���s!˪�Zt�������~J��,e���d6Ӎ�����	���Z��<�&䡼�ѭx���8�������aP<�TBb��-�m�k��`Y�2+�M�-'ڬ��hf��뢚9������@QPS�J�A�} ޸���}p�L_ys�i����h:�/�[]@T,����7�)���c���i>yS��p�����P�-�&��6%	��!8��!{YbL<+~�dm^�����p�R�� �29����XysH�DFd�]G�`�hCL�Q�=~� ���\e�|����z��J���~�r�2��v����p]l�3��b�p]���^�OIN�k�D?hUd:Js%��C�s��I(}�Sǘ$׌��n���m?8w�q�3�$3Hbo�A�UML���Q��h;b(�/J���*����R�цj8�FF�H����&���j��=���K��uV�nSsՖ����G��Ni���'�b�U0�x�y
�M�b��4 ����7���YŮuɫ;q�%�sZ�!X8�����t��e���#Ǆ���*J�ݒ� -�L���8��:;������I}P�ߐ6�C	�b�;�!����V��y��\�/� ��QO5����I����EFG9J��?��!>�X��+ꢸ��I��&�|#R@��n2*�@)-����"�&K�d��K�l����K��������}j���lޚ
C�1�?�z�Uk�zZ��*��3A�L*�����x*IOXLTZ#�Ѻ�aJ�@ma����qI�;wb^�t���|�k�Ї��CYm����N� ST�;�0�p��ыq��O ��p�C��������6�1(4Ԏ��0���b�u�q�����Gk\���]�[0D�����Kؗ�P�圡Vm�w�|u��O��Ģ��K��G�jD(|���zpk��é¨&���y���7D�XގJt��>�/l7���<(��1d/�����FQ�Fw�n0f�x�"�@<���{D���6s����O��53��I���W���#�V�Dw+b����i�i�Rb�0��S Z����A ���u
:䥨��#ݤ%5f�2�g7�w��͞�]�o0��怬�60ӻ���8� �efn��!,ѡ��+�{z��zW�Y�v%EB�C6)�]7P�1v�)
�6��{l1w�G*|��[r[Lx?�K�Ё$�dR����u���W�yX}��٦@��$�5��c[�0�F��b��X`���t�ɺ�W�9�=!�Xo�A�r\��3�bRAD���plq�8�L��E�PS���� �S�S9ڪ#�y-�]PH@��C@ՊўuY�/>�¦yʰ��"��@^�Ft��_D{���`S$��g��+,��;��j��,��DW�Y����}�S�kU>r�UuA0b����xƻ��ý<hE��M讛PR-*�$Z�C��T.rf��|v�櫜�}@�?�b����'#�!�c�ןC�<=��l�&����E�6�4�E�h˃�u�z�������E3��!��e*lw�sׄ�d|p��w�����&�S�� �B��j軔��RH5L���P��љ~`������_umy�
�F4��nk��|�/�#�\�eǒ\� �=����Ayf������f1��;"�5`~Q^a(m���c8=ۊ�"G�&>��b 	�"��g�Ƈsj����L#�~J�9
V����@�W�z�^P�cW7�p�s�U+�J�(�\���e��TѰ�8�Q��2��LS_N\%���d �f���0�I����t1�~tm95��M�Zj�!��T}k�%�Ź�bJI?�GH�J�#lX�Ǔΰ�ܕ��WZʂ^���nI3㾿و�f_'��TEz��0��,�q<��rQhn=U�Ti�S-��4,Z�_�������MLLE<��@���|	/�Ī��g���~�~Yu4�B� 奻}�u~�~;J
+�����G�|Wܵ<���h���ԑ�H�x2/��t#�FＣR�ؚ'ƞ�^�j?z�����Zg.n�9Z�E���+z����p��4��Y�V�1����)(3!����|f�$y�v��]j�iaэi{ ��Ԙ&�?N6O��
:�T��X��]l$�Ն���v�:U�KgB����B�?fm|�3h���⛞Ǻ�\@\2jcC��_n�����v�R̎����?">7��X�T8�2.������%%P)���_���Y@���BɈo�v�"�HFZ-ܔ~�A�=�==��I2k�:$��S��{)�:_[����i��Se^e+�wS7�.�eW���;���z;tb��k~S'i��	�k�N�p$���J�f�����z���,�_�q��M�I��%�'���4��"��d�׉]?�B\E���0�\��/�;-�g405f��d-�1�=W#%�V� ��N�16v�����i�Rn� lE���n�����R�&:���\���y��<,��l��]�V�X����;���$�������Z>;YkS�1���m�Oj� ���>L��\bV�i3��#]k�l�7�ǭ����j����s��� �"��oZ�����k�y�� X�,5R��q����+8�A���>s�ʳ}�YG�t~(�|D���r���Y�Ag�?&��ޛ(#�2�uie40O+���!i�3n�B#��(���z޾V�X�LYn���v���?6�z+N�H��NO鳾��QAK��t;���c�K�^*� � r>��yo^g7�=Y��	D�-�t��}l�ÑbS6����ly�a��$�Ok�5�AK�ݵ������k��V���+��t���M�$�0��`T�)��:�B.���R��gU���+M*�UX�V:��~��0���>-�	0M���Űw2k��[<�����>�_�Y�k��7�z�#5B2�t�?����A�:"!����V�ǜ��	X�?��}uC������+�x�jO�/q~W�$;�����Y R�kSZL!������>��@�T �љ�U�Br� �π����:�A�\�'H��RZ͹������*�+��u�� 9�-���1����v�%2.0�L�p���ږ�z��	�������%�_st�9��1����8���x(ۧ�zJ�8�t���96���fslO������L�M��|�.�3�Èr��V�+��~��<bʜ���[ј\���[{B{#~�'�<,�?�	��A/H%���~�VeB"훯Q�����-�M���-����l��r`F{IF�/F�`�����K�!�U���M�CUoj�������qGr��??�s'�X|���z���.UV*S�9��3�$�H0�*��Ҷ�Ӟ�rw���uG����Z�1Ba� ;�>�_�20��Q����7�/��1���Jv���N��&�v�1�����G�׈[��"�*��h�m�c��^J��T�:VS8l��^ZO�ovxؚmP[p���Z(B���A>Ÿ�Ʋ/�\�����W]�c���eL~��̙�BO�&/6��#M.��¹&�9Lû��=E��/�Z��3��G1�{���E!�y��Å1�����oܱ�s5�Otg��Tc&Iy�J�m�v3�o��]Ov�O������%1���~�Ov������O���vq�o�T������tBҎlϫG�E�+!:2�L/�����jA�;��x��Լ=����D'wD�%ة^{T�����Z�=^�α>��7��,��t����KzLÛ>m���&� �p�=���md��`�c���&+����W��Qs�^ɨ�0�&��۫�K�Rn0o��`�>wA���� Mw7��Vs���NR-;P�g���T����HU�H:(�(�W&r���g��̬HL=�Ȳ)��ךS�|�-��%}���X�x�(�3�7D2�^�q��i�^���,��E�k.�S֡*P|�R�]b�]F^lcL�O��Rر��/��|���/�	[����5���ֽ>�;��>22����f��#��5�oq���t6��<�S���A��O�i�t�i�~ �;a�j�R�n��?Gqk���`�;�PJ/ŗ�!?��Q��Y���6��D�aKYh�Vƹ��6���
��Ԯ먣�t�&�؏ԋ!�D��f
n�N��Z�?����[��^��+��$͕�t�# ȐPT��f��Ȳ������ RN���7߯P}o�:��꽇�m����<�T�{�;����C�,�p96�
s��<��r\Q�h:��	qr�מ)����e�dɻ,�-��ug���Х�kЇfמ��"�SF�(�������V��4'D,�<�sE)X��k���4"�]�5�D�6�ԗlZҶ
ѧ�W�(^{`B��o&�t��4 �BX<�Q�������TG�b���Y��קS�d�iY�4g��3���Xr�o����#`|����)V����^m��7�
n�]��=<.e��~������#N�4�U�L�G�l?uɊ��ܮ	�e��!�?�_f���'(I�f*�T��B;x&ԮG+<��Z�/<y#q��_��#���%��!�%�ᓥ��V�}�'7��(B 4�I@WƧ��}���UB��EQ�=����9�g�_8n m�X�z��e[c����)
�U2U��m��yf��"t� �O��\G�SA��q��x�BA#��!%��[����N�<a���;����Z���;��׶5=L��G�UE��$&[�Ӿ�q�*j��h���X^X�]�u3  d����bVҀvt�	L�����49�j?�Y������?��ox[����z��a�C!P�̨M��Y�h�7?-�`β��{�?j�� ��X�p��3J����#��0������{��6�0nuB���i�%>>�m�0"��g*����d��V4nwi�tt$�H[_,�?���A2��zT.�Z�ܰx=P�n���p��T��ŢU#j*&��<�y�d�&'��