��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�O�5t�"!�� �RY0�J���$��x�+�D9���m�P;\�<�"g�W�	x�k)*���uj~��H�wLj� m��I���%�k=}胄��<�v��J�޼1cS�h�~��X�?��PR%rs��8P�W��F ���-�R!��鷧+�7J��j�f�ͣ�H���5IT�������B��+���p�"W��j����4t����O[��:.u)�-�)�u~o�~\�y��Dbm[CN�愴Zל��<�S�Z%La+��<��2\�4�o��QU��� �cm	���K�u��/3��ٴ*���S�i�8+��m��\޼��`�NBBe��y9�n>,`�ّ���6��=a>$]����铺P����!��~��tq�|�σ��n�Y��"��p�u"p$�&L����sL=2<�{]%oF�B�^c����l(��`���_q0����j$��͠����X7�!�����Bq�.�7��Qx�Ԋ��W�(K���Lt�`�30��f=g��>33��
�2`3	�]t�:�KB$p&��8*�zkI|��+՞?L�ح�7�6�‼�ú���I��6�3�n*�鉹�C�n�Rw�����R��a
��!�o=�'^�n64�@5��Wi��cI@����D+�	���!��i�����1�@�F�Ē��:���X6��'s`ˁ�`��Y���K��w\�����<���Q�S?��ܧOΨ�@5�G�j5b�qv�a�o����2�0Z6�ʾ���x��$�h�UQ}�ە�M�q��<|puI�0 � ij��؂D$�1�=ES�H�� [��!Y�zW��X��T0� �~�s�%�_�j�wò�V^&����\G�x:{������Wa%,�K��}�4gGYEg��������Cz��˃�43��������٫!$��k���\�7��d^��_�O�2������Jv�x,I>�����2U��Vٰ�Kɩ0��?�����cx2�<���-#]!��Ni���w�A��2q�jH� �s�S��y���	�3�+�4��8NX�Ս�buJ�.��x�̒z��|�/j����Mˁ)��o[�DF�A�頁e�����V���Ҟ��)~� ��}��CR�RP�9Ę�z�BM���`L$�R9Ft���~/�$3�V%�$��������߮�ot��0,�����M�ءpdy�Y�
NW��'qU�aMk���i���Tz��0P����b &�y��z���`�+�[�җ�G�؜.%:�E!��-��m��R��(�Y!��'�@qqf�Yy����x��}Ү4-��7r�bV�&�>�T�#G���ڂ 2ݞ�}�fڭ��Όwc>�,�#�c'�{g//v>ڱer�T"��_t-!L�����8��@k(Ɓ����W�ד(j��G���1y�V�&�R��g�|&*����<�RAYedi�a���pf�E`�lQ�?��o���%���h�jGd*�#�n1������B�%]������Ӿ"ѿv����e���y�v����J�Bs���b�Fz8����>I��V��3��_<uⶩm/jV��"ʭR>k�iN�e>�u�j�y���S[l:�V����E�f�� �A8�Yr�<��6����vd�u:+���s�@��M���S�5��6"���uZ�{?$�,*�\�6}�,8��4����@a(�8j�uo��S�?};��/�����\'�� ����UAF�O.�,����%�o��i��}�p�ME'̦fj=�5A�\kC`|����u4r�h����	�
��j[�D[�ID�=c.�
���h�o ��N߁5+�G��2����T@~�F�$�C�V��z���ⅻ-e˗���Ε���r,n�5M��@��i���M��,�$ᆞ�9������p�I-�*�!��U#�?�΃�?执Z1�m�/�m!"�1də��FY��0p�̇���G���\JP����bȣ��~�
�I] ��>{�Cw�J���˲Zru/O&%$h:�]|.G��+^*󁈥��c�Z�Bm&s1v)���5�_�w�,µM0�z�p�>���z+���Ȱ{k�}ˏ���X���4�{���H,�;����1|&�"4�R��Fy��D$C(Ho�g���_PbWlg]����2�F� Jx�)9�8��j[78ũ�1yׁp�n�z��h�����VP��K_vj����;<�K=�ӷL��o:�	���9vZ$g$��^ת2'��%�cLB#E�-�;�ǬZb=�(el�ω���>� >b���k��E"�FTS"�J_�ZΖϯ)�L�wp2q�Y����6�j��H�W����\�.���ѝ��:��x?� �.�^
�#�P��ՙS+�	�r֣�Tj^J�r���)vD�a���D�"�QB��ϵ�<�x�.���%����W)��!#�|�n�sϳ2Hꐛ�~�dP�ͧ�2C%%�|�R�/hyy��L�_��[k��+^�à�TE�W���t z�����V�I\�p�':�x"8��">L;f��<��D/S��c��{�52��7W�0m�dq��\���%��h��[�zz<�g}]��v�[w~U{L�|��s�'�o��c�}Zb�;څW��O�F���6�	�9*��Y�k��gO(�ܘ�.��qO358�p�ģ)(px]!����2ܐ��|���X��O6	NvX���U�'�PJV|�uS�dXܕ7ͳEt>��3��IS	������ԍ�+1*��	8Z����U������P�����m��03ٕ�v�^1�x�`d4C��o'�k��8�4
A6��|f.��<����G0��'ĥK��sQ��Fa*j�]�z����vK)��pA������6R���;}�*��;�+� $�N��������	��q�����̳襕BI��4�����fk	tψ����j��"�{Ǵ�~;���0���P�-��3	�uC�o~�e���`��W�nSΉ��r������f?��ڦq� ��Ζ�΅�s�j��g��2uz㬠��Q�&n�)m�؃�r�6�s����,θ/R�#P���.�AQ�w�҈���F�y{Y�x�tA��th����J9K�NҙI��Szܰ�w��T���jjg�Q�Jj^���pY�F��ЏWWY�qD�{����TL�eA�b���~e$C�<Ř>�cy	�:����0�;'@'�Wi4'%5����Q��*ᚿߍ�ԎvId��aZz�m�	\�6�j��B� �I0xq�F�I;/ XI"C��3u�"E_D��A^B�߸}���T�Q��L��@�f�B�,5u��v��N]�3�Y,$D�-R�ɅalfU!�>q��ς��Q�P�+)H�0��A�)r�N!��FB<��{L8���9t��.⫇�F-r1���.R��<z��X�u��6�!��s����[z�iY�hKJ�k��	Bt�kE�$��*�$c�R1]$0 �ޅ���6"қ����6��c-ߊ��Lb�24��LŒ�$y��D2�3"L�Z�#qM�hI����u��"��v�\d!���K�Y�ۗ3��ξ��}�F�n�I�6�Z�t��~�k�K �����>9�=�քp�<��N!��~$B! M͛י�5�m�|`t��Ed7G H�p��j��RZr5�9V�w�Ty���Y��d�|�a^S�z�ۚ���Zv('�������H�@3�g�/�a6����RE	���K8K�đw-"��.v3/�~��e��ѻPz�z��
)��K"����^�~�O����4OU����p�5����s
�A���^�}�{���Yu�*�7�.B�.�]�|�2[o�Z�$RKE,��<�MD�ק��LM9��-���,����X{c_PCb��I&�\SY�І�5Ya+j*@�pH.*���I��k&8�� 
��]4Է����75D�Ӹt�����O_&'�������5��a.G`�P�F
��Go�0��|=�7e}-�\��<76C�x`$��U�"X]���a�#G3�W�{�ǵ��iEC�x�Ǒ�&#��5��������N1���{?�����쐞"N&=�p#+��avt�6O���7�av�<��0� Iř�n�HC}Jlj-���!�Ȉ�f�Z1S��{.�u��	z�#��l@5_������ѡ�I �RDY� �lV���!�v8j�?6����h#��Nթ�l����'H0Ex�d��ZL��[���t��ǣk�:�0g3��	���J�}�}�c��Rq�:φ���y([wm0�1qa�nyi"�4�������BƷ[�J�o�9E_�=B��d>ǉA����-�D4;Ə*��?�Y�Y)e2ʎ�]t<QJ��!R���1��(�����w���=���.�!��Lmr�54�
ܰBza�S�#iNi�xB�I&���W�6Y,�'�mJY�_�[���Z��}�t>�CśHi�Z/��<Md��^׹%9}~���̵6�O�c6���U�r�ܣ�����4%_�a�޳-��
�9[sе9Jh(]Y��A4�����Ԑ�3�-���j�1,���~����6�)�^��E�E|�+���{���^�-u��9���0�ʪ8U₾��{�v�m�&������د]�b�|]�k*>{Yn�;�ⳙ��Gpmщ��m� ��2}�߭�\�l���6c��Mt�Ƨ��\}Vrra�V냨�Xu�DHƮaJ�H.G�1���Vh����V��T8B��]�0�7�/(��g�6b�۠��F�J�tXY_�^����C�%зJ�96c�EFA1���?�N���Ǻ�Y{�fG�j�
5�.�1�޺�K�۫���,�$qwy��Ub�A��zb�˗o��{iV�<�����H��K!�ݼ�|"�[~窱�3���Nuy��Z?�DLP��.���=뤉U%L�k6I3��On76�0�]e@L4����|�Wk��&|�u!��u���z��g#R��P)�1���A�B��>'|���=�4Z���~eͮ�s�4%�DFf��H�a��k���$by�����U�R<����K��cUf�!�!V��GS�b��!lJ�|^�8�'4��a_��t�F{K�l�ǧ�����!~XgB�g:]zv�n�>3
btx�g����k'&7^x�;X��L��O�y=��A� ���0*8?�#p`�Go۟�,�/���Nr��}<z����u����1>����hNާAի݂�[<) ���	m�K~�䧖uP�U�ǭ��D�	)X���WA��_�����!]����]�H��Mgt�c���`��ÂuR�9Sf9�˅�,���#~�7^��V�:[��&�/��F�-GV��Vu|�c��f�DMVR8��죪�݉�?[|[zn���U�H����&�iKjC�s8ŋ���~��@$�J���Ųܟ�O��kȵ���Ʌ!�:cY���o��d��Qs��:��6t�Ē�ùYr~x�ԛbg��J`{G��]����+<�?�Yo�/��]�+��R���g�sq�6��-^���qD��O�5�G��@�]+���}(���ڠR��Za����0u�&Z������q�gʟ��N����xt��?�Y�7�#>Y�ӽ�#��7NV�I��vO�%~h�S�
.����c�����w���jxפ,ڎ�A��j�H;��!NW��3a����,��G�&�x��и��Ӗ������|�/)��{�8Ip]h)����X���{�����K5T(�����q������M�(�2(�^9�0TD�z�p�^��M!D����B$��>�fF�Bo�&�@!I�hiC<4�^YJ��6�Mܳ�s������8������	dٙ�n0ds#]z����@�UF�HM��qz��?=��������J�%^ōMV�%@'\�4t�Bf{O7�t�̕��Q��GoA>/�ց�#���Uۮ�e��@�0��y��Bkn�k�:|@�:�^ъ�C��JA�J��;�B�D,��m0iR�N�����~����O�jO��+�q�Tb#%r�ͮ$F>U>و.����s" ��Ή�_�ɝ�Y����Z�)��lÏ��b���%K�}���1��Dg��-�r~�}UF��ae4�>��盕��I+�(��[7�"/� ��H�E��!"�V`��^�	D�%��cݒ?E�A��^�"/炓�P��׋�S|�A�����:qM��i���D�1?�8t|�ڕ�7jq~c� �8v����U�D^��&�/K�|�k��7�ŗt�6:$qB�GaBK����x�uEA��|n�C��0�EΎv�@T�ۛ2lS~�����>�/A�ŋ-íT�t&h��Iu���,�J�g�t* 1���C��� 3�P�EK0�8�U��b�B���zg����Z2ЦȊ���v��e���*6ׇ���۴я���a �T�&�^&��M_?�9�����/H[�?���0�o8��<ɐq��7E��^�n��C�;/()lL�3Qv<ΒuB.�'F��/��&E]��\j,����N�|��Mz���p:\�3!Ь���� �E�ꔾ���*������d\�N�\�ղ��6�_H��/�u���{��qH��Z���N�C��$)2��{l�R������Ǹ����U��>�Ț	 Ů5x��:l_���}�?�K1\��S�È����A&/���Vr>i&��2D�D��Tu�xG��ik_��	ʓ��d}�ɒ�A@�*�Iy��F�O �`D���8����:5�x BV��J��|&y>�@۰��/���V�Wˡ'��e�FHQ	/���؏۱����̺��83�\��L3�RS��P6j"/���r�ޠ�-3{5��_+��F��F��m���?��~�(��૝o�VE�Ɗ���I����K��/>���g$�7l�@w��t��D���1>����`�j�l�k����o/�{��ǘ��Ս���R��.2�yb9�#gT��iiŀW3�_�n�TE���9���t�%*4lц^���ݧ�}Qjc=�$����If���)���9Q���ʑ<���jh��.���ji��$�B�2�����;Nf ��B���[(�?j"-t�إ�W��ZD&�,����VG%�n#@ϫ�#h��-#h6J|��j�Dʦ0�������
�)l�6�|-��X
�3L�I]p�#�W��@]���G��y���k��=V٦	��N����T�s�׶5Q��aB���i	��<�><���W�!3_%��*��?���m��$>����oA��C?[�￐������=�P�C��'�*�1x��a��|�Y%g��:�Yh����S!&��U�c]��[ե��K��JG�[��.�Aī@u3Ĵ>�����X�;������S�G-�A(��_�UV�&4R��(�(+�g
\���]B���m7��ƙ��;yͣW�?���	#�N���p��Z�<��1�_�}^�b>���~�n廋��2���d~�	T���$Z.��$V�8�}E��k�u8�����=��/����d�~��� dO!�{��]=aE=W0�
�H�e֐;t-֊��B��^H���n�[3��n��~N_c�e��1F�b�DM�Q�F���%b�o��x.�`��i��������[�W�`�Ŗj-�H5fT�n�U��
8z�ICX�Š��yVˋS�k����V���hf�_P�Pn�$@���/�+��ˏ����"Clr����D�l�Rq�� ��g:�)!!><���fӪ��w֏�����_�����K�����`����2�2�Oo���37��Zռ���U�m�W��\tDv~�ۗZ_���SZ�>�-ltOj1���sR�N0-9��b�#	(E�Ǵ��r��
[�<=�H�!��pd*&�>�X�h�`�-=�k��0��aEϾl�>2�ѿ�
�hm���W����.y��~*
5��n�l�Q������������R/��qp����9[Zñ���W�ٗ�H7Ox�o��Q���#�.�3�`����O�0�o�d�4	���d�Rsx�}CE�]������t��ֿwά���FQ�S2�KU����7e���i�',1��;����J+���)� ���."���cl.мB�N��v��=���7����+��
 읃|?���\_Q���IY2;�-���O�EZ-�6Β䅃��{;pó������B�vZ��Iڐط��0�t0���b�������,�ӥ�E	$����syy0����:)�pm��|v����H.��J�:3�s�V�i�'O���3m0�9��┌�8 \A��u�#ck�?�(&�W�6��}Lsn�}�aR#ś��ˮ�٢q�4����[P�ʴ�@�t�8���,����ܜ��`՞��al�0�FZP���8;��:�DrH�<-� �e*�49�.I�]s�~���H�=�yg�h��׫���B^h���`��ߦ���(�<�\U�l�'���?��`�=�F57M���y<0�Ai!� >s���Mo����,^�,h]0 l��:�#�XcdѫSaz�� p�;'���Ď֌;�����2������
�����҇���W��X�UPf�����uz}&��d�Fj
*̢M�ZA��Ո3��B�/ɓ���ϡ��;�Zz����q�9�vx�T�g5Jz5e�<��	�i��S��~��i�Y����g�:2�p
x,�a���Uvo���(��@�\Eĳ� h��$��������J��t� �h�AC����Kx���P�w�!�a�$_�t�ܻRNP��-��ː���@����*���d��[Ljp�x���c�������$��\�&�r�I�*N���l$cܙB���D������/?���yZ�r��6nV�N��!@\m1>�;�y����8ܗ/�E���������`%��UA�vM��2�w��q�O}&]$T��ʧ���l���x��8o�Y���-⛲��V`�t�� ���r�`�c�m���J2&�Hҷ�r�)�B{*#���N�a2c�-W�W�k�����'zAm�5³>�h��w����\�(3v);��z��	w����+L*z�yj�=)�oe�O e���XY�����h���!��@z�߄fO��k�^�|�$��3��|v#}�0��u�`��u�̶I���d��@��T*sS!�h����_��pj.��g*����!
uP���ƛ�q��M[����jcӸ�MRYJ�{8�F�$�����N=ǖ��������q)�K[o�zwr����3'1���`y��e�&7�=[:�/&/C��D/�*��ޅH�i?�p����g"��4m\J-g�Q4��U�R|���"��3|�ѿ�#�Jl)�!��	:��.#��LJ��GE���'�//(qN1�
0�1q��>�`�%��<�G��k��8����I���_�]+�'Fe�&�:�xf��}_�t�雬7i����nho��^;�����^�ϓ[kz_�~���������?����5"�+��
;��ۺ<xd��j��Wѳ��h7�H�Jlq+�t�%����j�l$r�Te:�r-+��AabH�X��w�#�Q���r��.�*��$\ �v�EtP���L`S��%�efv,*�˛ �7�'�W#�E���4�j
1���jw+���T���]i�����};�'�qb޼^��j��:�1�B�_.U�4�j��m�G@�R)X���2��m#�P	0��=��_n'��;R�����b�$�|��"v��	v�a��`����J�V�Q`��4*8�%��%��FL�/�������(��L^���Ҫ�lOx��&�
�K���k]���Ed�ݣ��%�]y�CU�4������3�a���T��ф�΢�N��l?��SB �:X(����Ws
\쥳�����/��x��X�yƴ���y�w�ߤfE��AKܫ�7�R�'��(M�4,d#4�w|LO�����E�E:�'�AVE�C��.Aɓ����jml���X�a��\�eA93�u]��hX�eKՙ0��)r�_a��[����f<��/T(E�K�'��hj;��x�Q��}W��J���g ����N��q���<.��ľ-�0��ۈv��9`Xݽ\���d��O �n����E�gU�\:�~n"�Uӗ��2��f��|8���&�g��3BO��^��Ǯ"Y�i��~�b���_!@��B$ǫ�:�~�{�b�Dǟnz������`�#~v�Oa����`#׵İ@�7F��o?��pO4�<ߜ0�l�>/��ОJ����a�����۟�01I9&����YP�6�u#�H�ɶ�W���+l�k�W�2Ě&;"���[
�����k�M<^�ƛ��(�����sb�m8�!){�T�P��E�� �#��D�n���/rr+���0՛v�X,�	�Ѐ����$�dr*<O��6�/�����V�L�#fc�p��%��J~ݕq��}	s��O� h
CD�_�_���������to9���M���E/
�N�>Jw��0������B�̱"vr�����ً��l�βHq��
X�����W4�7tl&1��V�]9Kl�8�n�M{aUE&�Ƌ\�o����s�����r��A��+U�nixΘ�N%�^�_�r��PY��O���X�l���;z_��3��!*($�>�}V�%ED��&?��G�#~}1b�W~L�q��Y���$�/�U��0ȣ֙L���Q�a����?MBIL^�~������4�ޕ��=���=H��{އ���Tg9������p���u&��~>{Q�!;����B��k���I�s�S1c>4����s��_yN�%��y����I:��@���9��%R٨	歮���ɯJ.��6��Y������C�|�\�V?hZ?�uI�`�rh��-�S��]O�%s_�x"�5s�m�L𢁛����R�Ո����E�V� H%\�n?S����n-	]̔���U��Za�:��T��xܝ�N���ߍ6��"����FEO5�H�?+���$��ب%�S_�=M������I�� %K�G Ui�
U}��V��	��#�SW6<�-?�)�Hʤ)�i��/��Yׁ��Q� ��/��Ҟ�̺�^5J�zX���ȹ�"��7s\$Γ�_��Z���FqlU��q�0{�F2�jf7u��DQeH�Jj�ya����-�V�),�H&g����[/(J���2�-k��:ru�D#ݪ��r�*<�Q� A�N7�X���)��ƀ�:?J �(koX���_��;�%�R?)�Z���6q�ͪ����ߋ�HU]R�ca��T�B�@�9���t�G})x��d�h�����ڛ\?��U�q���j����)���7���$�b=�~re���Ý�������Y�4�@���3c'u&��Ld�ж&���m�Է�'WA�7���L'q�I�p�};(�ط/e��8mP5����h>}ʅH�����7�1zX�j(�.��P�9t@Pؙ�FN����6f�>�NW�Mͥw�|�@�M�D3r�F��/����b��������%��sVj���KA�6��(�i�,�W�����3��g�
�-8Y__�������8�5��v��1�I��=�a�6��A�Q8.Ų~�\~b�y��'�:�k����l od���\��Ə&���-�]�xU#���s₭|�Q.�Ą#t�7��p5V9�̉�%O�˩v��]��E�Z8-���9�#���ge���y���,�}�[�Tݿ}Z��'���(cΧ�?! �h��^����j���f���T�^�=f\��O�[����bE�m���d�^�/U4�8b��S�%z���H�6N�̥�_��S�M6��@��h�N+������ij: F[&�`��c�F	�e��}c�1�w����)ۅ�Rd���ƚ8��k2�Z5�p]p{�|�j��S�>�̓0�<��f��s���B���>�w�=����%�/�?����h[��������f��� 4�#�Z���q�g��!����OhM���w�u���Ǥ����{�����K�Y��C��U;{�~��굨ԈI�Y������\e�p���{w�x� $`N_�c����#�1�'|eLH��i�+�^Z�O�}�����l�2$�#�M���0a��7�7��o �Vz�a��M3Pq����p��ܧ������Ŕ��_�_BB�8.��䤹�gA�۔�%�
W%�v���n�dUख़s�>D��}�������se��4�6_���Ę���X���L�p^����� �y<�^/���R+�I����P���#x�-�L���1/�)c��
�����>	��;����� ٧������z{` �d��s'����ǄRL���Y�[i����4i=]{f~YZ;۝0��sh����vS���,[�Z<�r�(P5+��M��y���^g��?6+��sy�L�tC���\�h�W9�>�Ep!ø�u�}w�W���ИJ��������X!KL�#�S��|��B�����ۢ#��l�%�2>���)KI��3��3��4��4Tk�{'͋�i�Я��t��`��-Pl�'i�R���:;A�Tv,���&���2����d��#��wD���X+�#�8��7 ծ���,�����Ω�lC=A��a�o�hB�xA��ڜ�ʓ����22Ҏ~RD��������_=PC4"��q�f`�%�NQ����fA*"�w��|r����"rm����(fC$72+���t���Ҭ��֬����QL��}u箵�K�T�u��i�؃��CJ�6����l��#W����^1���Y�|�� �11-Mo�E�<�p����������i�� ����4�8�ZM��$%O ��|��B��@��+a���Xx$o��<�U�y|��o�����:0YS>s� �9��:B�$���5V�q}g�dM@��Qa1}C�"�[CN6�}���_��)�@��ֶ>��� 47h�tQ�7XpΚG��	� ���iP
B~� t�S+�!đ �}�qd׋���w���H��O���	�QgyCA�ܺ�e���9gQ���a��%p ���&lyt�� 璒��*n_�[85%;��i���̱�YE_���cr���?v��_��dX[G�JqÒ�w��d|��W82�=��3"�({p]@��[�Vn����r�4�9�2 ��sͅ��c� �I!B )*�����hh"��=��nR�7�v�E3 �æy#�+T�B�Ŏ���F8�A��5��x�x��S	@ye[ǧ�S٧�kpѿ~�5k��,O:��@�NW���òD�C�rߢ���J5dG(�n���y����(��b��Jϛv�N���Zl]
o��~��@�92�d�^�[(J�:7�3��"�ɹK��f{������rF�\|��w�O�QEShC9�4fI����MW��.�H�h驺���Z�EsJTWe�l1�a��_&�~]A{���D&�7��I�3jlt*��y�I$@��O�n}��'��gGwg�������h\f�B~FH8�,%���"n�T�ep�lFƮ�R؏�1�*��Bt�^��_�/�T��%1�1��lW@�G�`Þ��$CEѝ��2;�r��R,�Fp���hzw i2���z�����f4���1��Rr�#�K����h�["r���+�Lr��
�.U��D����7]�Һ�%�T���gU�B�_t�� ����6-��j���&�x͖����	OH`�E���8�p�1�������c+���ҥfJ��f�o��52���_V�c<I���j!���)|^�(t��ּ���~�&K�r�Un��W����'0�?*��Ҏ"U��Ǌ��Sz�|����1�|�J�[/\�K��f��#�CqM���!�y���Xv-�${[�������n�گ�&!��]�#�n�2�߉��`�f�~���������<a�+ ����®[�ME�Ndp(�`��"C:P�e�$��H����0Ux���a��7"�kLI��kv�>Jh-���^y-uX>^v���q������Ҙ���Q�ɸ�g�\wĵ��z���hu�?�Sng&X>�B� ���f�2���o�KH5�L}/�
���K��!�(��a�4���Ξ�2�~���~��tM3c�#v�,W����m�F�Jʖ X�=�F�o*�=��O���_�`�3��Q��qs��c���W@q07��c��K=�`~�c����o�����\�o�"UB�I�~�f&:f�T�x���~�,�v�g��Nq Z_�~���Yu��ӇZ����L�DL�Z�y1���V�ϋ\O���Mx�� ~�����h�A[�7�u*�����?�w�Z)|��1k�T��h/".��E׏��).���~a	�R�ϓ'�C�N�o܁��Yr M���>n%��o9ĸ�l �{JN��D|�d~+	���h���[��g�;���g�!�^%A���S<9���Ƒ�����,��Ր] 6�$a8�<��\�B�.�j��c�-f�U�2�p�{�9�b�R��Y_�NĬ1����0y��Xj���c]�L��)pîl�F&L ��f���4쏃�!��5��:���.�c����I^���i��%�G1���|R��O���Kh��S���ջ1=o���%'Z�Qb�t^j]�ǽږ�Y(�;�_�<�D�O�>k��*ĳ�H�@�!��>]���M�3����pA<et��rk��{��@��:B=	j�F�~"��+% �$R���!������7�.s���Н�7��w��v�D%~�mn��8���S�t�[�\�k�V�t�3_@�\QJ��o�R�nA����0~~��)��S���Z	f��F����J/R���%v�{;w|8��o�C�y�uE����M���*;�O�Kɬz�$���3`�y}<�*��$(�6���.��Ox9(k�_&���ѵ���8d���L`���3�:<1����m���7�E&Qg�:�~�jDȞ��YG�)I��.�#���Z �;x�Cv'�B����\1�bI�eAF���\Qd_�,>����A��C.����2��e����	�����b�/��~�ڎ��+�gT�����Qy9m�h�qX�u���������Ո�:�aea���f��=3�(֢z���'u��}�]Z�fkܹ
�q�R�u���n��#�j��O�
]"=7Zz�B/�ǜL�{羶�`G��O�^,Uj��G���<b����72��%~�(�C����Ϡ�T��x�k���Y��Q�qF��$��u��l��~�®bw!N�, [j�q�L�U�V�[lڣ��$�_W>���i�<��݉@$�;�v((�d垵��d?.����jL��(��GvD�3+Sæ�;�OJV���j�X��@o��b!�`֙qH�g�� �5ʊf�k�<���ɛ��
��n����ŻS���l7p �1����f����p5�^�u,.țS�����+�=�A ͇�cX�4/Cd���,kzm��H�t6����{���õz���B��sE�qp�V��\<ނAj�β�y$*�e�8#��E�������c�q�JX ��R�^�w�uv���c���D�y'�
�)_���vsɐ�_��yT�+lƦ��y�6-b⓹4M2׫B�͚b��9�T� �Z�'����&��[��u�����l΁�J~�������������uO��%��/��bDp�#_Rj0<�%*X��\�s���<��k��ѝ���L�vh��Q�!R!LW	�S��p��}]1tV��:��;�46�Đ$z�`t�V�K�!:C����
�E(�\�U���T��%n�i	hfl	�C�5�@��UT^E��=��mO�W;=�sH,i x�6�<�4��M}�-�b����ӛ�)}h+1�՛�ΙZ�.-�XI�kǅ���@^��{�L�%���O�ڣ�B?.?��'%ͧy�E¢A�;�q���!W��Vik���C��m]@������l��%D��U{~�{/ϣ������O��Zpr$9���&�1tU5-C�l�Q�!���I|� _"܎��=��'��V;�=�1�	��Y���q`��˘j��*����<���ql2��$�P�k^LF>�	��Z��p���&«sYE�9����l�ӵ��&-�z����:�z
`m�^��./�8疴���Ek��=�8�i�.GVd_?�:�G cģ�q�<��3`�'󑊅��t40�̫���.k,bA��⪥u�Ad�ʢ�s��?đ������ �ղĕץi\h=̡�#觩3� ���""[uս���t|PH��nO4��[�hx�s�Լ:G
&[���K9,zxW��@O( �D��� ψ$h�����$q[۹�-�>��26q��_jɿ����_�l^;G=`��x��VIMAY��i�1s±ֱ��"6�x��;RW��f>^B������ �A1נ��3=�T\�[��Ղ�^���Y�:�467���TF(gO�5{��R�������.�yjA,F�3�}��4,��ւ@���H�?�/����di^AY�]��v5y�lyU��/���RyJ�y��^1��?�����RϠ��UE���wV����>�K�Tm@>�G���b�$^^1�J3\ O�O*{bͦɀ�]�����4޷��!�8ܸ�q��-�0����D��b֦0�|�J�������;HB�qqkg���a���4B��2 #�!���NgE.N�L�9�p�dZ�3�������s9#Y��b`�����U�����+)�z�ZQv�n��G�m�QJ��m��"?��ܒ��Q^�ġc��U�B�'*#�[i6.�8��3x*zw9X�Pځu��v6��&l�IU��<�Fl��?�����=��BjWeL�0�ǘd�,�~Υ���$����`�v�=D�Z�o9zY'8�V\��*�gp��H��,І�BK��g�����$��P�h_|y�0�E'�o+�����`.9�e�^$f�nN����\~/K���?)٠B�1\���o��[vWv�{m_]�-��(������VuwLv����㏀��ୈTw3�qq3��P�q��0:{k������oAHs�y�ҵt�χ�v2}*9ߵQ�O�&�1����R�)"�z����R��B��䜟��->8�­�� �NQ'����&���g�W���6l�����"��,�o(��F-Wʕ2�7R�����b��W[�!OI/���XJ��w�@1yO�����m[.\C�J1�!�m[����A�U�sRH��k������|U�x�$����E��W��Z��>�M����7e8�$J���f�u/��H3��hUs��u��ȇÂ���_�f�����럫F��=��y:�)�lPͰ�>K�1ls���6q�w��X��5�SN���d��g\H�)��f���U޷a���,k��i�&��/�H�_֞ah�� 8�5��N+�����+:?h�~����,?��J�!��G��}"-fm�ȿ"�(XL�E��C�q�7�E��� ��B>i��L-�l�IG��4��Mm��ɤu�p��QA�Q�fˮ��'�)����R�@d�7�˺u����`�u�6��:�,\��Q�\c�z�o p1r�Z��j}�0Q����y��z-~��h��@30���
R����|����� ��$��o&H7�r����ҸuܸF��j[��ӫ�|��]�".k'0"�ֺB;��(�S8
�^�~?X��a�D�'�;D��������Y�KID�n2�������Q�9�۳�~m�Q:x�׾��HD�2��6���Ɔ\�v�6C.�xLq(Q5��,>Ҩ��a�H�m�s��n>Y�4-e��Y�%��kR�@+b��L_H���R�ZV�"S^��g�"p\��͍^	�(ZkM�l �#+d)��k�2�dJZ��`�}��y0�	���qnJX��lr��O�'��~���}h�u�Z�n��s�ɸ���4TE^���P\^d�3z֢޵���d�CT���}�����t�q<A\.*��@��l6@�
�Yç�}��,�,s"q~�7��`���Ȏ���IR�^�O���]#�M,b���73��p�ʐy*UIܼy��Ql����'D]CQ��w��D@S �2��߁۽��)�M��K�DV�w.�t��B�M�F�M�G��+�h~���8s",�-T��PQ�C�Q�g�"h�8�:���kc�xa���c����ǯ�Ex�_#C萮YN�5f�0��F<z����u�>5�Zѩ�?�r��%M�)0�:-�Jq�c1��ĻF�W�}��n�L�e�"���s%%\�<��y��ґ��"к.~GK$-v�-)��㊃k?R�ב.��LE!Ş�!rFA���Z'�3��ا�*������0�5L��#���+�P�n۱K��
/��_��;�寏>Jd��)mm��
͐	2�:B�c"��8�!�ԧ��8��ܓؐ�mĨ�}�%���]�٠�mW}���r�d����We�G�0��F��S�T�V&qԔ�0mY�74f����q��e���$�7�őX�2�ئ�⁝�F�uT�:đn��$���Ж������y"�1ڄ���
߆��A�R����,�����t�9�Ly�H0V|�����T!9��qc�K�|�Ö5\P%�%�� v��P�^(�d����Zދ&����2�Ų��#����q\Ž7i�?x��5������ό�k��8�S}��U)�ɮ��黷u�2N�V7x؝_�tބ���%A-�<*�8S�u�	��U1����J�^%ʱ!��o&ֻ������ �f�f�����S�[_�X~+_�
�E�;"���V��d��W������q{&!F|�՞��Q�LkޞOgj�7.�b�Q|]L�f^���lj����	8G;��Y<�;��{ӛ,!�R�҆l+�Bc��nyԧ
/2�$qޠ�<:f̹(b������K�/�N~���1.�ꋃ�Ȫ�e��J�z�2"�2��b�����(-�aQ��*�L�dfeD��)R�O�~�i��sAҢR�;�PwJ�*�^ë���D�Syz��~��w�X����:�	=~�c f(^�f�%N�����>��R����tGio��!��Pa�%�8�mΑA+��������'G}�s�� �Hu�A������b��bv�-xڬ:���.)���]R���R2����U�� �>4 C�oi�lx��E�ʹ��D�w�C%lm��h�z�/'��	ǫ��|��Rg�lW�d鉰AT�T�[S<]��%iQ�ב?���JB�w C�L1ځ��	��'�+�Ҡ�����53����0�]����?����Ţ�۔$��ڙ���g� D�7~��D��>�B�*�Qe�Ϗ���:�6$;�0��ZG���)Ӌ&_e�r�E댵��]D$�Y�ˡ�p�շ�dFʷn�Mz�cĄ���U��%O{�2
�N�f���D��K�B�90Ȃ����^����s�B�ɽ�Q�$����.�΂Z���Un��מ^[3��0�n��*e�ü劭\�Gۏ��N;S^�a� �����
�kZ����^ǭ����0�cI��&C	�%L����K���#����@������F�|� j�+S%&Ԙ�hx��쟊�nX�N�s �Ǟ��i�����*���w$k���]{��)uil� N,�F*D�����אx�ӵO���YA☂�D���a2V�f\��ZV��}\����Yp��3�Cu�1ꓱ4��b�KF����F,����4�N��N2$���=�3��x��v�uL��-b�tTdAoiе��<��{���7����Ԗ}�ڝ�T�ݡ V���u����R��v1Վ�f8����|�Ruy1�4�*|�(1�؏�H�Zt�~�6}�>=뗸�Y��8SdR嘫���4� Wj����B`�79%_̓�(�v4[B�j�o��c%9���:�j�K=��a!5C�-Hhd*��s!��y�����(z͡)��4�� [S�Z.,��#S�)dc���m�co�= rr].JB�-���K��:)z�����
�p��*��c���pR�?g��B*�&��ڙ�4�G��&��E���xÌǘ������`� '�XN����09�0���6 �<P#��lNu9.Y���G�T2�ϯҾh�w���2���Q��U�K�_$��gw�~�Jԓ�:J7�?��7�YQez�s���L����3�m�KG,@�A_׃/!���]�0�^�=TR�G�ܗ�G���Gwm�!* �C��Tl>�����z-��t�L����9Н�@�5������h,w�j.W�W2��� V�t���{WV��p<��K����ȵ;Ϸx���{�**���`�D=A�we��_֙qj1}��GUKO)����[�jW-�8H��Fr �k����P ��1 �\f���
�I遻5��S���JA/�qnm��a���4�$��EO䍬tnׅ�8k.�QuΏ%�>�HU�o�< o&~�E�TXG�����܅�<j5;վ�����ِ�����#\%�u�_(W�F<�%V宵9��z�e��*7a������q�i��оtͭ�nj�M�2��eZ9T]ҍ����)��~H�M�)���%�������v�;	��-�� rkH���:p
;e$"��m��￶����q_@{��`���P��rK,��=�!Ʀ*��iقT�Og.���J$�*\���x(��DN�nm�FV���<�8ʈ�W�1�4�v�=Ɉ*��k8ts�`2��ܽ���ܱ@4��ŲE
L�1��e�b���MQi<s����XvOn�N�({�.��OS�L�SG#-��1�S�v��Zc}s�ix1��֠IY�PK�-i����J`�w,�J/�@Ls����t4v �"욠�a!4.�@NFhfBSل4��N?J�2�K�SI�)�^A8���#Մ�ﭥ�]��l�<�z۲�����o��]�n�e�]��������c����_��m��)V����a�u��h����h�DVn�f��l%:ǥ�9��<���� �+�9 CjQ*$}s1_�T��\�߹���;b4}�%C갥���~�G<eKy��lC�9�dڙ��1�:qw�'�qy�,�Bg�fM��Y�J�Y�:,�ը�afqL"���@���9E�1�F�]�����v(����T�dZKW\�|�i���~�-��G�*W� ob���*���&q��R؜U>����0�Iwu�B�y�evPQ}t�B���Iэߪ�������Lg��(�a�},q�"3���7���zI5�Q�瘇�Y��l)+���g����-vӋ�Z�J�L+k��c�F�fq�s���
�~��湎p�#��a��z��b��s����"ђ󭼗�+�ж�գ�s���
q�'��H��rj#'�HҊ�&���/�'0)sqK��j���%z(��ωp����l�1�2{�u�ٍ��ּ!�П��9��F�k�wE�"�?IR�666�һ��呕�����2�L������7m|A(9��^�:q�[e�b�L	S��"L3�ۜ��}v!�b�r'�O�?[[�����w���:6���S�'1����qL]l�B�z��S,הr_L>r����e�]�K\ąV g�L�x������`G� �A|K\�y;�����D{��z!�LMá�V�/M�[`xL���D����u����u1�(�/oţV�(K�My��`�T��E�����c����/����߳��B��z��g��R�f�*�CKw��}/�����2�T�Y�#�؍9�l��XB`�%�T��dƀM����=�LC��e�A�x��Po�-�Y1*Z��D�c�#�ʼ��8�\o jC�(�L�k������� T�b�����ʟ
�`��L�����D��4%��"V��\�����:ŃS0ւOӇC[}yvfP�U�َ��8��1N�Y��?}�)�!��e��&�BH�M+�|��ݙ�"��#j�0����cP�|a�?�w��mt ���!�k/ި��
O·��vr��R��%�)Mqd�p3/e�r�v ��X�-���e�����I!Si���'QR>�pQ!_*(+֧���Ƚ��#���p�Wk@��S+ʺ����E� ��{�	��VU�>�
��v�'8�6TċMH�OY����W�ϽS�������,X��ws&9��zR11
�2#���.�� ����2���m���ۢ}ե9Om�<���u��6Os�[���D��S����lj�;㉅Ur=v������7���e�IG�|��j�K���>�f��C�.�*����n��~��Q��L�RW-�~E��̉i7�{�hH�F9�IUb�PQ�����$����t�[���U4�d��C����a�IC�i��o���ݴh���%@���Zd���m��a�?�����lǊ`#��;���k�^��u7�wtCî4�-�4Uw����:dӬ&�e��ҭ��N����؟D��@�9 t?��1HyZ
M���N 4�<��"e\ T�Ŭ����dI�c�������p��
�D6msH)$�).���Cw�a�&���-����ߊA�+V��Θ# u�6���G�'M����bQ�sN�z�X"Ow����|��<U��\ت�έ��y�XKcǫ^N��	g��"Gqm��7nm���N�\�j����ڠ?݅?�}�q���b)H%�O�f�c
	��͝\\?˾�+��n��,�f��7O���0����}�|����B�U��UL�V