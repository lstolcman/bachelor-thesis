��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J�-�4ϼA�IŠ��#�U�(�f���+�p-Hv"�-L��wUoV�5�󷹿1��4��[c��i�>�cű�A��&;"��+p���N�'�p��gMG��6l�7ֲ@eo2;��5��_<\zڪ:C�EwZ��6�&x��Lq?��n]�9⪎�o�PE�G�k�ڑ�O��f�;�̍Y"�)ߞ�m̷����#.��؜)�	NY=j��R��#o(��2W{���,Z	�H��Qkٝ1���0p����XR!ξ��,R���@��@���E�BcF�V�K�����`>ol�cAG����{�Zt/g�$�e-��KL���nW�ᅋ���hbu����u��7��\��@W���7�7?���22�ϵ��a͘�hXR�^�A�\x`�K���`��/�i4*+%��ʽ�w}��w��n����m���d���5=%���G��+k�)��qK5��@*���$��2����x"�0+ƍ�L��-rc��V�(��/K���~�M�a��{���ZCҍљs���.ս�����gЄ�y�7`�`w�G�����P_!�l͜�-yG��[嗅4��B���i��5�j���HL��W��C!8�u�T��޿Q��tB�cސ�	�� K�9"A/��ru7�2�.ݍ��M��A=�"R��u�< ���1�)ᤢK�l|�ptA8}v���w��������'=0�DŶ�����3�0 7\��� )�!@ M��j�����v�������Qg.�v�$h�M�w���(H�S2*&O�����ͯ���,���_���ս�z�����"\ ��:Ղ�e�	$�9#�츪v��������)�7Te��a���r��g�?	��i����X�]#�O�?��A��A�Z�th���������&.�l�w��� i6��$�&�+;	-[{\!�$�U.Snv*D��I��(팚� 8*���#�M�p��fV�PaˮF�u�<������o\F���-eKdE 16�z��m����-i1��b����[�'2�G�ϳj.��-��ND�U�����C��"��`�'�,�mpQ�������4F5�OE�*-���kI5y�#k� u��944������x��`��!�ʣXX�!h�F��i�6�E�E�hj~��)2yq���f���p�,lz�.3��ZƼyx_���,�{���z��J�2��߱QV]\�㋕�e�(H� ��NfL��s&�I���1_���<.��TU4��������6����_A�J��4��q�!O��uRJ�w:��P��7�uĠ�{[����	�p:�"7��!��-f�3lu�wX�t���@�������Q(�]��ɦ	��.�R*y��uR�tH$���k�2M��H�W��ے$8�+ui�S������8��;S%J1	��24�;��"�M'0"���+X�ѡ̄�ch7�g���Yw �,1������k��B8��w�����̆\Ñ�[ƐH�;c�|�"��z�).��i�r�UN�Jе�������^c9Y���s���lx�'y)1@X��]*wӃ�s.f���DL��$}�_<�i��i�����@�Ê�"N!�<ΐ[��!��}0M��s8�Dv�~<O���9|��/���HY}����i�ƍ��w5f�ғ�h7d�X	xt��犯��x�� ���g��� �����p�����-��0KH�x�f��"p�H.��%H��Y�83��ޟ�S�B4k8I��UtEo i*=m����L5aQ�BQ��7��z$S��\#��,w�<�x�b��P�����_̲t(3];�.��sf�[�c�V��l�g�����軴E�r'K�&M�äu@}	R�)�d�='W���[v�=&w���b�n�6���|+������	��Nk,I �q�K��P��7�{|�Ly���FK;K�LZ���-��T��>�)�e�"n�U�� h���g�nxn���w��d~V��V#Ց����c����Χ�QR�md_[�y���J#&�}t�%��I�ca)6�O�~��X���ɫJ=��3�M�7��o�7��Ek�pw%}�`u���;����-*�8q��A]2 i?�,m%E&��yw�E�� n>�Xۛ)�'83�G��Nc}���j��G�����.g�eȁ�L� ��Ҏ�ݝ�F�>h���n��������ޫi@ת#��#������.%g�K�5�ߛ�sl: � ��w�F�~仾���$�B{?f�+�H荎K+��'��s1�+;��>�%�8���1^ΐ�5��ӥ����<ܹ/ސys��f���/��R�n9��=����w�\r���U���z�*�~����f;m
���L���6]�,LT�o�ʒ�bgܧl�*�}o%���`��3�����g�(h�U
�=Y��b$��c����C��c*<d��n3*_R({}�sp�=g��7��_�3ڠ�u�U�b�k8z<��:��]�%nK�v@(��NF	�w��V�����!����\N�z�J��ge|1`���=�V�U���5��fԜy�����y�����MD�����޾a� P��)i�^�S���Dk�_}?X�Ե��^Nh������!8Q�.(��Z�w������G<��c�l0u�̇��1���!�:㰩�O0����ޠ��
;�[��F
VEy�����Y��aj�|��ze�(Ŀ2
"?v�-�{sM�t�K������q������IU�9��țgܰy�X�����`I��1�8\���iԹ����PB�(j4���U�F��&	OV�t��Q0
�F=�j6�c,�cvG���SdS3)9(�?SW{Ǫ6������O��C�=;��gZ��^���p�ǯA�N��!��T�	r�ŗ�o	Ψ`�? �R]��%�'�)�BLm.UZ��������X���2���SB��6�0
ݕ^C�.��j�F%�lS�#��JHӥ'����C-�$�N��/�xz�F&�>64��Wh����i��*:y2�_7�3ִ*m_ȞUڶ1�zQ)�Y=frw�a=�||c4Z��30J��vv�����<;�򝷄�dd�dv�3�SE"���W:L�Y���CW\#��F�N��z�7~w�8^�#�<$�u���I:&@r@�G��������e��^��ʜ�� ��a��}ǃ���1���Y@���K�Y%�c������y����V`����VZ����>3� ���mbrv=4;����p��?�|�H���Z
�Ǘ�4�:��^D;˫�c�,���[vQ0<�n���%�5w8�`�b��j���945��,�O��:����q�U4�26e�z��帴�D�mJo�ɉ�7Y�������Cu��{�����!J�`^�
h5H�)K���t�`]CڧT�Lt"6ʄ߃h�~xe@��
�_j|x#��7�pcPz���&q��j"Z�u�Y�jߵB���٫�,-�����3*��E�:�z�f3%KM+�d�E<��"Pu�QϏ}:�V��|���-Z2����1i���x]9ad��BjM��W�h{䩫h�cP��n.��[�^2��{�����p�.:�[�OS� �b���\�:*�iz�@J���,��ĭ�KS5��^�M�[BR6�{A�5;R<RKK�m�aN�t5!����u@�.*�T��X=|���)<oV����"�8���j#>�$V�ch�Q� M������WL`;����q+������B;�EB�ei���M#!GX5�ɼ�'W���}�W@|S����S�l��y��3��sn �Ya�İ��̑�5'=b��cLу��GWv#�)4�x���0���5s�� ��(j��Tw[��ʂz��h�Wc��]���A����T�K�\�vN�����Jx4T�W���GF�|��k��|;E(c�>� /���$���D���b�vӺ���k>�TaE�k�9-K=R�	��Ȣ��7
�	��'�[�S�9�����,��b�|����fc�˞"�D��8	w|x��f�&��@��df�ȁU*��kZxN0�� iԫ�@a5~��Z�ڣ�>��,+V,0������38�2���N⸫R����4���	T�v��/w��B�������<������iIO�V��,��8Us^A�J�j]^&�mo�i�9Ŗe�u�O%���x��/`çԂOu���Xsb��4�/2&�������=�z5� ��z�,_�B��p���Fd�64�j�c_��6�0��j��7�q��E+��H�<-�9�1����x����C��*��i�$�
_����xM~cI��sP�e\����z�_BU^�+"`�0D/M%�R��eK�~���Fj�XW(�9/����㝉�h0�ȑ{p�ۉ��<g��@�r˸};)�$S���u���a����M`��������@�w}b�����ɜ��N�.�f.��%'mi�D����%7�Y��^0l�

5��k���p��:F[�#��208�<��o�0������|ww&:�U�ܛ��'�F��~(��c*�=׌7~��)��5f�'�䨷m�^���������7�+ĭ����u��P��?���s���Bw�w�
݄��p"o��?�� ^!��b�v�\v��%�nY�K�ʖ(���)�����-�(�����a�13�	�uiC��&��~��I�5(_�	�q;���2��[���j1���t�H�C�]1�}M�&W��+�DS�@'��C��:-�=�mqq���ƙ(�7�	�v[ P|���Y�h�Rn�:.��B��.�S����C�^%�.�L�w�z�1`S�
p�tC:�{��#��kR%�6�l���'����.���;�r�+�a�>��p�I�uN��8�U[��②��aa{��	݂n�&��WG�?��U�a�*BE��0'�O��:������ZA�\���D�)�Z.�c�p��֕�Њ�{>Y�,(Ti<���s��&P�y��m�Y�یS|���#�����/�4/!���µr���S�1�Q_
�����W!�+χ@˚�����P>4W\���1eh����V��?��;��Aˬ��x�1�Ed�&��k��U�UN#yX3�'�6�"D��l������'����Z ����'�Uk5F�T|dUo��23�M�{ˁ���(�]Q0�1i���]ŵ��V3>;~�@�h�xp��ľ�Λajr�
���$���_���W�-�~a�bBG�*ּ%��$��
{ox�[��`�i�Z�.c�ǰ#Bh�2 h�������!R�zս����b��>$snG@�fY�cƙk�� T��5'Z��u5��}���+K�$��޿cL��������I`�~���?���1bȝ�s�!�k~�/���4)b�qCA��[3�Kg