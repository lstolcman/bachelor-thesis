// megafunction wizard: %FIR II v15.1%
// GENERATION: XML
// fir_first.v

// Generated using ACDS version 15.1 185

`timescale 1 ps / 1 ps
module fir_first (
		input  wire        clk,              //                     clk.clk
		input  wire        reset_n,          //                     rst.reset_n
		input  wire [15:0] ast_sink_data,    //   avalon_streaming_sink.data
		input  wire        ast_sink_valid,   //                        .valid
		input  wire [1:0]  ast_sink_error,   //                        .error
		output wire [22:0] ast_source_data,  // avalon_streaming_source.data
		output wire        ast_source_valid, //                        .valid
		output wire [1:0]  ast_source_error  //                        .error
	);

	fir_first_0002 fir_first_inst (
		.clk              (clk),              //                     clk.clk
		.reset_n          (reset_n),          //                     rst.reset_n
		.ast_sink_data    (ast_sink_data),    //   avalon_streaming_sink.data
		.ast_sink_valid   (ast_sink_valid),   //                        .valid
		.ast_sink_error   (ast_sink_error),   //                        .error
		.ast_source_data  (ast_source_data),  // avalon_streaming_source.data
		.ast_source_valid (ast_source_valid), //                        .valid
		.ast_source_error (ast_source_error)  //                        .error
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2016 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_fir_compiler_ii" version="15.1" >
// Retrieval info: 	<generic name="filterType" value="decim" />
// Retrieval info: 	<generic name="interpFactor" value="1" />
// Retrieval info: 	<generic name="decimFactor" value="100" />
// Retrieval info: 	<generic name="symmetryMode" value="sym" />
// Retrieval info: 	<generic name="L_bandsFilter" value="1" />
// Retrieval info: 	<generic name="inputChannelNum" value="1" />
// Retrieval info: 	<generic name="clockRate" value="130" />
// Retrieval info: 	<generic name="clockSlack" value="0" />
// Retrieval info: 	<generic name="inputRate" value="130" />
// Retrieval info: 	<generic name="coeffReload" value="false" />
// Retrieval info: 	<generic name="baseAddress" value="0" />
// Retrieval info: 	<generic name="readWriteMode" value="read_write" />
// Retrieval info: 	<generic name="backPressure" value="false" />
// Retrieval info: 	<generic name="deviceFamily" value="Cyclone IV E" />
// Retrieval info: 	<generic name="speedGrade" value="fast" />
// Retrieval info: 	<generic name="delayRAMBlockThreshold" value="20" />
// Retrieval info: 	<generic name="dualMemDistRAMThreshold" value="1280" />
// Retrieval info: 	<generic name="mRAMThreshold" value="1000000" />
// Retrieval info: 	<generic name="hardMultiplierThreshold" value="-1" />
// Retrieval info: 	<generic name="reconfigurable" value="false" />
// Retrieval info: 	<generic name="num_modes" value="2" />
// Retrieval info: 	<generic name="reconfigurable_list" value="0" />
// Retrieval info: 	<generic name="MODE_STRING" value="None Set" />
// Retrieval info: 	<generic name="channelModes" value="0,1,2,3" />
// Retrieval info: 	<generic name="inputType" value="int" />
// Retrieval info: 	<generic name="inputBitWidth" value="16" />
// Retrieval info: 	<generic name="inputFracBitWidth" value="0" />
// Retrieval info: 	<generic name="coeffSetRealValue" value="1.38088023046E-4,1.57979655075E-4,1.79163289322E-4,2.01675075698E-4,2.25550539965E-4,2.50824509531E-4,2.77531038845E-4,3.05703334529E-4,3.35373680387E-4,3.66573362433E-4,3.9933259407E-4,4.33680441576E-4,4.69644750031E-4,5.07252069848E-4,5.46527584035E-4,5.87495036355E-4,6.30176660517E-4,6.7459311056E-4,7.20763392573E-4,7.68704797891E-4,8.18432837935E-4,8.69961180812E-4,9.23301589851E-4,9.7846386419E-4,0.00103545578157,0.00109428304348,0.00115494922276,0.00121745571381,0.00128180168557,0.00134798403731,0.00141599735746,0.00148583388545,0.00155748347687,0.00163093357188,0.001706169167,0.00178317279054,0.00186192448151,0.00194240177227,0.00202457967497,0.00210843067182,0.00219392470923,0.00228102919598,0.00236970900535,0.00245992648135,0.00255164144906,0.0026448112291,0.0027393906562,0.00283533210204,0.00293258550219,0.00303109838726,0.00313081591827,0.00323168092606,0.00333363395497,0.0034366133105,0.00354055511115,0.00364539334417,0.00375105992532,0.00385748476254,0.00396459582342,0.00407231920642,0.00418057921575,0.00428929843982,0.00439839783319,0.0045077968018,0.0046174132915,0.0047271638797,0.00483696387,0.00494672738965,0.00505636748975,0.00516579624804,0.00527492487404,0.00538366381652,0.00549192287299,0.00559961130115,0.00570663793211,0.00581291128509,0.00591833968366,0.00602283137299,0.00612629463833,0.00622863792411,0.00632976995384,0.0064295998503,0.00652803725611,0.00662499245418,0.00672037648813,0.00681410128228,0.00690607976108,0.00699622596775,0.00708445518204,0.00717068403668,0.00725483063259,0.00733681465246,0.00741655747256,0.00749398227268,0.00756901414377,0.00764158019347,0.00771160964887,0.00777903395684,0.00784378688128,0.00790580459746,0.0079650257831,0.00802139170612,0.00807484630885,0.00812533628859,0.00817281117435,0.00821722339968,0.00825852837136,0.00829668453398,0.00833165343015,0.00836339975633,0.00839189141411,0.00841709955694,0.00843899863212,0.00845756641804,0.00847278405659,0.00848463608071,0.00849311043695,0.00849819850312,0.00849989510083,0.00849819850312,0.00849311043695,0.00848463608071,0.00847278405659,0.00845756641804,0.00843899863212,0.00841709955694,0.00839189141411,0.00836339975633,0.00833165343015,0.00829668453398,0.00825852837136,0.00821722339968,0.00817281117435,0.00812533628859,0.00807484630885,0.00802139170612,0.0079650257831,0.00790580459746,0.00784378688128,0.00777903395684,0.00771160964887,0.00764158019347,0.00756901414377,0.00749398227268,0.00741655747256,0.00733681465246,0.00725483063259,0.00717068403668,0.00708445518204,0.00699622596775,0.00690607976108,0.00681410128228,0.00672037648813,0.00662499245418,0.00652803725611,0.0064295998503,0.00632976995384,0.00622863792411,0.00612629463833,0.00602283137299,0.00591833968366,0.00581291128509,0.00570663793211,0.00559961130115,0.00549192287299,0.00538366381652,0.00527492487404,0.00516579624804,0.00505636748975,0.00494672738965,0.00483696387,0.0047271638797,0.0046174132915,0.0045077968018,0.00439839783319,0.00428929843982,0.00418057921575,0.00407231920642,0.00396459582342,0.00385748476254,0.00375105992532,0.00364539334417,0.00354055511115,0.0034366133105,0.00333363395497,0.00323168092606,0.00313081591827,0.00303109838726,0.00293258550219,0.00283533210204,0.0027393906562,0.0026448112291,0.00255164144906,0.00245992648135,0.00236970900535,0.00228102919598,0.00219392470923,0.00210843067182,0.00202457967497,0.00194240177227,0.00186192448151,0.00178317279054,0.001706169167,0.00163093357188,0.00155748347687,0.00148583388545,0.00141599735746,0.00134798403731,0.00128180168557,0.00121745571381,0.00115494922276,0.00109428304348,0.00103545578157,9.7846386419E-4,9.23301589851E-4,8.69961180812E-4,8.18432837935E-4,7.68704797891E-4,7.20763392573E-4,6.7459311056E-4,6.30176660517E-4,5.87495036355E-4,5.46527584035E-4,5.07252069848E-4,4.69644750031E-4,4.33680441576E-4,3.9933259407E-4,3.66573362433E-4,3.35373680387E-4,3.05703334529E-4,2.77531038845E-4,2.50824509531E-4,2.25550539965E-4,2.01675075698E-4,1.79163289322E-4,1.57979655075E-4,1.38088023046E-4" />
// Retrieval info: 	<generic name="coeffScaling" value="auto" />
// Retrieval info: 	<generic name="coeffType" value="int" />
// Retrieval info: 	<generic name="coeffBitWidth" value="8" />
// Retrieval info: 	<generic name="coeffFracBitWidth" value="1" />
// Retrieval info: 	<generic name="outType" value="int" />
// Retrieval info: 	<generic name="outMSBRound" value="sat" />
// Retrieval info: 	<generic name="outMsbBitRem" value="5" />
// Retrieval info: 	<generic name="outLSBRound" value="round" />
// Retrieval info: 	<generic name="outLsbBitRem" value="4" />
// Retrieval info: 	<generic name="bankCount" value="1" />
// Retrieval info: 	<generic name="bankDisplay" value="0" />
// Retrieval info: </instance>
// IPFS_FILES : fir_first.vo
// RELATED_FILES: fir_first.v, dspba_library_package.vhd, dspba_library.vhd, auk_dspip_math_pkg_hpfir.vhd, auk_dspip_lib_pkg_hpfir.vhd, auk_dspip_avalon_streaming_controller_hpfir.vhd, auk_dspip_avalon_streaming_sink_hpfir.vhd, auk_dspip_avalon_streaming_source_hpfir.vhd, auk_dspip_roundsat_hpfir.vhd, altera_avalon_sc_fifo.v, fir_first_0002_rtl.vhd, fir_first_0002_ast.vhd, fir_first_0002.vhd
