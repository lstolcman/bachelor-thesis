��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6��Mg9��X����6���
n��U-"n�ϋ9�	K����Ӱ��k�a�MN'��d�D����%q8��v�+�dc
�"O�c��R%`��Pt4
S�����}z]�0n�U�Ni���+�!QF����~�������J.9]y��R��&|�Ή"w��4ф{3؁Z	V�l��R/Q��ւ������D��5�IA:`��~y3�cf��s�
%��Hy����}�R�#DĈ�c�ܿ�͵O���+^?Sv�M��4�85��H�DT,���"�^wOT��vB��rV;��LH�	A�S�����)�b.VtKXؚ{~w+��s�PI����,�$"���D���	Jĩg[�Am��r$\���x:C�p���u&ȼ������9d$+�tu�6h'�?�m?'	Rd%Y������Y�-.���lYi�]�}t��x]4kd�~c�R��v���!�h�s}HA�R-G��U��'���������������ݫ���
��=:|�'��
��mįV�!�i�h���
����N�nm%3����e1'?����9^�)YY:��B�6�maE��&/��BK� �X��+�٫��0��۶�Yu�I3=�t�u��a�-����][v˺��2����˚�ZD��<ξ���3Wq�B%�|V���l�NF6��E��Ow�&�+�(#�d�����x@�>��`bޟ��ɷE�4Wf5�eo�B[��V���٭LwW��W�.v#��B�+�B�uS���֯��3in��#��"��j��Qs�F���ˊG�}�v��D�F۷�v)?�Fpy.�w��4�����B���Eu(�`���O�ԖV����<��1-Tk\/E���"uy�M��O~��y̧�}���2$|2[�����&�=�ӥ�n1��9)�9��}��B,���v�GNj�&�cj�"�Fe~D@��(�T�>�deb>=����Ք�0�~&�f�l7�|8�^I�s����w�NK ��䮗����m�~t5����2��k� F�!��-\|%ҩ����8���®���'��-|
o<n�@ D�+�6�(\���j�1�M���4�=eL��L���J���^��Y�k_�3/�@�q�Q_��Y>���4� CX�����:3밺��6�g"�Nu�`�qM�~���6�����lt���0$�ÕT�ڑ5
�7 ���r����Z4MK鹩?ky��|G�D�AFP���qF��[H�ǛT��rE*��\�g��`R��k�������(�K\&V� $�ȇ� ��eo�	�f`'�t [	'S��L'(��XQqc�j��<�3�kD#���cy�.�
�8�]�'��f�����<�Vņ��?������ܜ�=���߀]��QTWӠQm����>Ӝ�`� �Ӗ<n����
�_eL�ld���*��w]vc�Z*3-�f�?�U5���x�(rr����Y/gM1�U���,'��10'�ەL����{��O����M�ǥ*/�:��xy|\���CODr8�dz�X� ��/�CM{�L��B�����ڋ�XA&P�����ȋI�� ���~j��]
�W�ɫ�Xoirp�V�u�VaOmT�$��S�.���,��D��dy�$2%n�H�mG�H ��M�tWZ�33ٺ/;Z��	�m��Ԁy������(��2�����k<�����6܅�������\EY�h�Ј:LD!q�*�r�0$��m-67�Ѽ�<�=Ϳ�0p0;��C�̷t��Ɵ��஀��d��0*���������G,ͣ����ϛ��q�+Gk�?67/b�@���b��O�cv�ƚ��~�&�ŏba�۷����s܌V�����c�h~�@%�ҕ�?�&��>%@�/�����}0ړ�lv�-��ͱڑAo�qF��1>g�o5��C��r8l�Z�ެ�Q�P�ķ�e�_�N{�ώp�>9�s��ꔂ(��h�����M�wD�Cu��,�?k`y�OY)}� ����_�*�FъI}2�ֽ�($G�#}x�G�F��$��\��RL�o+a�M�w	~-:ٖ�@�FO�r��=j�_K�'�g
�V �ֽi���KX��-W�id�6?��<%p�au�|�&.'����J���P!e���N/��@ygI��+��Ϣ��{?	�ʻƚ���,��ӾG1i�����}/f]�à��)�SJ(�pg6:n͆���c�jKTH��� ����H��h'�r��DΊ:��-�Wm?i��8�P���
�1���1t��S���;}$����>?��,�k���Vr�Z���A���B�އjB�v2�5�*����[/�p�G�ߠ�x�:�� ���6TQN[z�R�=G�s+|	ɔc�X��$�tc"?��g���l�ML��L��I*u7���ᄝ�y$�ej$s�	]��1���ƕX�OU���)�E
��k�w�pgG��dۅ��SAE�>;�{��xx|g4��˭@�+`)&��Pq�(�7���|� ���c��k!2�����#Pw
�iu�[7����A�ʼaV��3�lץ���o���{�Y�-�I�Q�P�?�����f�oܒ1�X�=�bO���_+�pO��2  _�3X�(`Y��B������G��Kc���E�l��wC٘�_����}E~�*�W�+�qJ%AV
@�4#��#����2��#6�u^���`r�(�[��f՚�G$j���W���`
��l2�X�x\�>ȃ�H�)<4=�}ࢫ�"|P��<qp�0��Bݣ���/<م*Xrh�WsM~�쓭	��Xo\������ݜ�X�-�L]�Z���Zi�N���{ы��"rc�<���Ѥ����Ő˜Z��L�&�:<��F^�s+Hx�&�Cf]Cܖ��'d;�WG�f=��$͜��l�R;�gk�ͤ���_�FEZ��#�j�=C�"��*m�A�])�q+Bj�6�a�x�r-�h���V�f�Xk��ԊB�y�����r��+��,w¥�@�B���dV@�?��J�-�>JkJ��4s/L,�M�L4�|,9%*�˯�+bAP�����Ӄ�ޏքm��Z��Ԟ��g.�a��%����b�!8�;�h��u6�������OKĉ]$�Sec����>��<��W��^�L�pa�LV�8�(����B*�9h�9��I\hux�S8t�
Q��a@�3ںX�`���~��R%�ě�U�Xa3�q�}z�<eJ���"b��WE�F��m�/��P=Jz�ǎµqM�R���s��RX%�����ߞ|�^����>��?pa�h5:��p7��1��m]/���, »��+o4BՍ�U}�:�ι�h�����><�D@nn��v�V������z���F�_΍����׫���8���}��/y��s��h5��M�g;�l�ZA�w��#�\{|�N�i�NZ#)w���SE���7�L�0w��.?����j�Aʰ�H)+G�|� u֒���^���7Ͷ�kչ�]L1a�F�u!���A|M9�`�:��9Ϻ��O���m�e&{^VM�3i,#��6V�8r�	�Y���:�����y?�ڃ�W�j�'�GA�hQ�7C�@rn�)O�܇�붓j�� �
�\0^����P.���5@� �p �a�̳|%!P���k���`���Y�|�7���	�ӛ��ݼ���x�{eD?Bm�^��ą�^�TJyy<+���ۖz�͛kL�VX�~�v�l�ȅR=#�C)��m��3O�Na@7đR	����>%��E(��˸!Y~�=�� ��@�R�($-4t�ӄ��K-������nn +����Ol��8�������4~��WN�ȩf#2�K�=A�4���1T�^	k��Tny���L�i�� W/4�2>�G6�V�H^��jE������H����$�=WQ��Ѡ�xA	!����Õ��j�]���3���u��o�"�7On�����}N �8���E�*��&l��NW3[���Cx]̫����He,��Sb�u�h��dC��*ZA�<� h;o�{G��e8�Sx�������L�n��40�e`%� �)pw�`��0܌7�'j�.A���=�����uε�ё��ڻfI�XU��f�`[A.��"#����Y1r�D���+�则�A#��BX�+�1z�[����mA(}�� �h�.�����V3��Zy��G������Æ��=���	���^ F>�1�kF��}�m���".�E����ˌj�q�͌�鵞��(���ai渠�k�dy$��3')����BY���b�_E\���>�)eԌ����vP�Q��X�^޶��i�E��u	�P�ґ"VO"U03��C�6�+a-�����g�;�K΀f���ԓ~�?���K�*SW80Sw�Ardƹ�H�[����p1P�l�	����ci����AR�ޓ�yj!a�(Gh�c�U(>Uz+���ҫ�v"S|���-��7m6�'� �F�]�dT�`�����s��vC7F`<�=���P2��݋澋1��/�ȏ��M{���Q'x��Hy}�,�gR��AONQ�x�Ԛ��0Fh4���ko�7X'm����hb%Tg�+�Uig���R-�#{A�.�����}�E�?����rC��,5o\Jt[5�M��!qW��]����0Z>4N� �l�q����kdZg �*�/�½NDSo��K�A\b��;�@EЪ�3
���lc�E�9!�}�M%=���q�a�� ���s��&8:���@��S�*:
�*�(��y��:�r���F�.�p�!iY-��?旞P_�\3V:�z��#��K>����*W���\�%tJͭb A��K0��&�HM���z�WHܗ�ʒiRHK�8��?/o%gѬ���Ť�,h�.���g����j�1���G`�l�x��ܽ6ԋtY!��j�'bz. ��%yq�	���6?@i��b��j���$��bzU�;;�TrIm�U`*�S�n����@��Ӈ��X�y9٬�"?y��ڜ�wJ����J����Z"���������e]�q������.��_U�G�<���r�y-��o�!�4X�Z��^��1[�V"/�Xj�cZ+B�;����"���|������c�J�@�
o���fP��@��L�1��3�C�n��u�E,wSs�O��^A(��W�C`�Ⓓ��Y��6a�����AC��Q���?�+*9\`�����H����R&�HC�)�Nq5����V�(%SQ;_xu����	���7�&gz)�,�
x`��CZ�6���φ	4�R.����뽗��T�ٮTl�P�����ۧ|x1E͌������Sa�i�ï��������k	��c�d�����5�u�E��c��+={���NE��2@�n�n�\�}��~}Zcj�bm��Qk%kJa��(�!���wv\g�M�6"����A�u���Y�)���RL�J-�])�	咲���v�Y�ӳ���Ͱ���>F�
���K6ؽ-���Z��z5�P�8�fE�02���(����6Mһ��������G��c��U?�֙Q>h_�湒���؜<�_�ٙ�;U}�8��lv�	�X?�)�Eo��A�R���_�+�r���u~y�}���b�Z雈������$ S5�\�
W�lG��Xq%������)/����
:�(q��V��C�,�)-ђ�3g� v��v�-���~���_1V���R�2'�)a3���.m� ?�uY~_���x�J���[օMَ�vF�<�����zbS�S�x���R��Ѭ@�_q-�|�=G�̎a8G���>��kp�2����d�*M�uϓ�y�Lg�:�N�B2�w�����kBp�B�*�$������5"�7͠)h:�X�?^�Q_И�e�:=b!�|�����z���%?!�{�]�^֫گ�����X��+#7�J��r�j|6��m�����ɍ��Ă�{�p�X��f���ۿ�Z,(�����J��}��*���=RNq!ќ����)���F� {N>�����D��lf���6���X�
��\�?,l��=~!@���<�D3�*�~M*�g�;s�
&�
���O��q�Q:re\�5�3��:�j�h,��C��N�dK�Lq��i�w�*l*F:p�%x�<�V͍.T���㏺�2,�;�p�񪌻�'8�\�OuՒm�}o{HY絳���X,_���e}^-��мn@طEJ�>$NZ��L��@@�ǵs����YGޭ��~(�c+#;*����#�r�?&��D��w���ဧ�.��՝Zտ��k��������?ur��D��=_���%�`���T���W�[�j*a%���^�y4å��J�X��!��J�
4���E���b_�g7�u�0��L�2�z����O��[�Y�m:�S�'���SѸaM��Nm�QV���W5Y��L��үf��F0����Z��G���n���)�T�8��(Ǡu#�0X�ӹ�@�a�]XR40�������u(侄ǿO�R�{;,�.���1��
0'�S(9�2�i�+����,?�	{w��U���4Ue��&��d'^��^�YGF�D
����f���Hv9Z20�/!;c�5��ɤ��=p�;�����ԋ�|�M+���8c�<�2�Ȫ1�Ȇ�(D6 /��طzF�����@L'䮔H�������C�\l��q2Z�U�!�|H�'�ze�W3��t�8�ղc?4fz�_��;*�� 4Z%4�\R7����a���ed��(Jᵵ��7����:������Y�����g9q�Q
��΢;�Ҫ"GU!'{x�!A3@��
��r�����=�F΢#(W2����>��K�ygl��d�j�M��u����FΓxG�$����\��O�a3���*%�eⳉ�%^8ɟa���qbo��	�dPA@])\|H=dI+�_��y}&A�BI����&Y�x���7�+9]Ǭ�� ��/�~�K[vx9ݎ�M%bQ��ZƢ�];4�RO�#��d��8�û;�fRA@�a6^ \a���h�X�֔���-���4���
DЅª�*��\�ڵ6�m���-�O�k*�x�;P�	9Ͽ��ἆ�ۂ)l�
�q�y�4f�cM�����"�
H0����kl��Һ*�@e8	`9 ,��*E�,�=9�����VQ�A�(�;����S
����N&$�b�6��@34�r��$�g�D��_�Z+g�����Ɋ��Ȼԕ"��7�ٝ-_�W�>Pz8�6y��}���ɹ�@g�;̜h��{qB0E�`t���]�fyId�'��&������p�������8q�^�ㅵ�P��W�2{l?vI�{!e��P�6�ϟ �R(��)��f�o�����C~�ե}#E�2�!0"�qsW�F
"<�N�]<�R΂�T�c�Q%�oQ��>��k��1��L#�~��MW����,�1M[��i�8�����\w^YG��($���Gǋ�������_�!ju��t��dkX���E�ݟ;�?#Y;�٨l~SФDx�tV!ߦe��%k�"_��[��o�%�ø~%@��>�ck��?_�Ы�W�������;��&�[K�NP=����\����E%v������'a,��7ڌ�w���x
�`�eL�8�[�������F�?��Cm�H?yƫr����g�t~G��	�=esg�X��j�������$�0C��!��w�{m)LɌ��ֵ7��|��h�E��!�?(ך	e��������Q�m����L��-���$�MOP[
6�cu��4�b����!�i���|���ء>��Jn���nm���֝{YR�b���b�ء�L�;C�2���C�,�k� �r��o���3���58������F��!��nuJbA��D*Q�C�"o��2�$e,+4����A�~������z��HK6i�������J�P	�h��nYZ�&W�����`�
''bݖ�2(S叀�[�T(���1��H`�u��W��>M��83L�T��N�����h����)n&x朒�S2���z��'��������5��_��3�@AGE{�!3�]�9�©Ɨ�?MzA>�+��&�f�VXr -%ԗ{��E]�M�F_,�%Ɋ��%'��T�\�1R�h��7��F� ZK�pZ�|IƩ�r�
����3�_��菱CS��|�h�nO����+������A����䍭ވ���=*��^p����┟�p�z�`J���o}4�<���~����«
nv��L���O��i7vt��=�!	���޳c�*�*М��r��ɋ�\��\����ތ�vyBa��z>`Lt����C�;��u�ԋ��5ŽvP M[T�׸[����)3�A�rHt~�P����%ǧ]}��V�|�XE�R�I����[��܀��'��6���Ҿf���ka&���� �n6�O�w��J�%�KڍZ8���r���v�"����M���
Ͼ�Y�H�<�$q���B�̒[^B��8eR���5� i|2;�̸,�"՞a�c�`	���b~^}�U�������1�S~,ƌX:5M�|�-.����6���H�C���yg���e�Ӵ)��aNf�cT�}rA�r$֢�5���vC��Ѡ�f���5�����! Ԝ��Q�W�8�|KW3�Y!U�2��!�<�.іN�&1�S��F�$G�KI�\�E��A�*�gL<Ohs��#�8d?-���uA�}i�FF�
�|��HN82�p'��H���$T��Y�4�"S^�>4MV&�V��u�o��?Ȗ�W��	k�Y����� !�q�)h���0�f�d���CN��r����rk��& }����2���е>�ѥ��H�,��;���Mfg0���[��y$�E��g�v�2�)�F��� �7e�+����%��:L�k��G���v�}t]{}-�S�G�(x���=B�<_��^1��8
���o�^�k�=�_ܳ����<��sL.5�|k.��>}�B�'�&�/����:����Ց��ΰ�@��8����D�	�����D�s�%S�-����A�`̫�T��R��㹄C�d�P�%����hʄ���<;�_�2�x{K
}3t���4�}3p=��Z�7H\f�94>>7������M��l�/1V5� a��00o,���m�����t�r�b.8�!�]�����n�L�?����!>u!��rK=�7���x��(bg���q,����	Al 8PY�[��d��(�=߉��(�Q�V �6f��ac����_	iuK`���x8!�m�q�����&��u��j����54��p������Q/�9��ers'�0hJWxDՊ }���sS�Q���a��b�}~�;b!go;�;����@=B|)~���d��� v�/�Pǀ���R��>e}7v��b�A��,�/�[ֳO�ؽ���{~r'��Bs�r?֖�CY#��1��]�v[Wx������r6��u'h�4(��3܊�4d�H\�܋+~�8��P��[EHÐ;CC�{10�50�׬|���	 ��_D[a�=]�RS�Q;�&��.{��lq]�]ரx�0Ga,2(jg+���_��ce#঴ivGi�A��F�i�m���X�<
��@�WE�&��T �P�3wX�8H��'vv���)!܊�6�rwG�&/�
���,W�-�f���|ݜ�̼X��RJm��F��*��E�6㨚�q:#&7�����E,�Bt̂�2n�\�T�/�(^�o7�[!�锷�R>��p��_at�<�H�Q�<'��W���N`���C�}����0��9���ťA�2�)�`){PՏ_�Yr�7}��m��U��7�"��s֟z"�r������H}~ ٠�
ܱ�	ʤ�m��R�ş��O�vE��ƒr�|G�}�>�&���o�Av�*=�Q=�@3X�y�ˮE��ڶ����2�+I�g@�Z�4{�@��@�J�o��d���^�=�p�l�"P�2��Zrtvz��?!��l�x���������D���H=0���~�b�����P�\v�Y�Z*�t(p��{~�*��{�󶻝�U'@9}CērH��2cdz?��T�
�A�r
#�L��C�թ߀Z/a�v�;��X��ߚ�\�x�9�\U��'���L�0>vM#�ӓ�w]�d�������@�-V��H:PRD�u�@�W
P,nm�p�Ke/$���c=��~�qQ���Rk)F�`�{v�ݾ��}�����vw!�����W��n}��U��2N��S�@Yq�P3W���%(LL#L�1�SZ�f��� ����R@�NE���:�ˇ�i/2�����p�*�lQ�"��͈bh���.fA� ��E�&��1��+��~w����R/�9D���^���(�&���Q/L�Z��R���1_��<��A��(�#c��B��k��[g�X�q�M�0�B���z�t{�<�@n5�M�}�9V?��wv�L�8n�mY�Y��c�9��H���`'L�zPhLڽ	s�Z.4�^��Bĥ�e-�ܣE��R^zT?>����瘤TӖ��Lk��Ɨ�bn]�ue�cyO����;�$���+.^8���?x�o%w�o/�4؍ū��x�r_��D鈨B�-C�|���
)Ļ*6)IfѼ�O�YFc��;:w�L@,��yР�@63!�n���:�p2$�&��#��|�JFW_��uJf��=&��2f��Y|N �f��а��ٓ�����q�cg?�oc�@\�1Z�t�%����b��:h��i�^�PXϒH�?�f}A����Jd����A[9��S�gT��+��������l���������I�oڬxjb�b����B6U�Ƚρή�އ��8�R��/y�Cnͣ���v��(�A���b�P�c���������.M�� �7�� s�	CU^NE�^��S�P1��Q���ؤ���^����k�#�T��[s�rR݄�H?A�M��������P}4Sℸ|�ޓU��L"�������k��G/TA,�#F�bDm �z�œ��Js��!P���f���cY��c��]:�)b����Z��E�7�~�h�}�Di{[kk8/
��'x}S�1"x�J��F�ǆTʫ3C?��_h��IO�{���ۏ�]hI��W��������~�yp�Y�R�x�8x��!��LhN��p I^ޒ�Vq?l #����;%��K�0�H`(+�w�V�Q�Y��k��=x6!�֮6x�q�������X����L2�r�_F�h�Ӥ�צ��#&
�� ��hYv�?\O�v���
ve�7��^���A�����ۑİ���'or���)��4\��'����gg���DJ<�Ri�N�Gd���#xr����c�4��E5�_�%��*X�(�d9*P#��=�G�O^���N���":ީh�(�c�*�����:Z���)�N�Gs�h�����#�"��W�z˕��d5�?%�O�ۢu�-�8s����j��!|s!8�hg��EB���>�ϵ�2���gfΜ�	W0 '�+��c�
wj�Y��r��5��gP�y��t@ Q�z:@��f���#N�=���'�u�((埕b��x&&!خ`<w�tm�1H��y�*.zf��-9r5�%��L�|kt���+�g����QX���:�ed`8;�08�&����2�W�m[�,Ȳ��R���~�xA�����Ҁ�
[˵+/�v�_��5b[�hFY���A���<���q�Db�3"Ft��2� ����P������* 5~��{�<�{���\�7O�/rNˋ���1z�1'@re!��|�;M`�;O���wơ��? A�嘰�S-�����Z�+����~����$צ~K8&@$^�WՉ@}jNUŰ�v�(P��s���&���͹�5�,}
nE�� l�n&���ؕe�M~aF3�� ���rʸxd�����w��G!s�?W�S�k�������A��f8�婯ұ��t��~;�-�h�ݱj��n8D�W���9���`�[��ߤN��~�4���A��W�d��X���R}�5�4��k00)�����6��u-ώ.����ɥK��b��R�*� ��5��|�+VY.l�CO��"���p����p[|�����]5H]�/J�<~{����I�����0�J>��qgQZC����q�%I���t�4+�'�2��c��s�٪?����"#��n���&2Mz���r��H'��[=$���9��%ߖK�!�P�z��q�fL}p�|B�R;�,����k"�L;�w��k�l��!+��P�jO4�3����t楾��c�%��I�*kg�2��L#A-K�NZ,h��P�Pr��y(�Y��l��Y���U_�h3Kg*�jN�9��ľ����x{Vm/�bY�6A=��$��щ m�@S��]	9"��?ӓ�4x�hy���ꇰW	��L�TA�5�ѯ/+�,�Qe3��U3EG��^��Aпv���ό~j��x��O�O�ܿ;�ߦ�M����U��[����ĵHSxA�b{�sMF�;m�
��
'tӷ��l��a�/�[r4"+�=Sn;���`Yw敊�B�}�g�l�`��+��6�������:E!�i׷j�n��6+ZP�6� 6��>��)rr�kf�;��?��O�V���7ӫ��!�rs��xna0�yuT'@t�/[�It%�ˇO׎�%�\�ڛL�׏���T���}�څfk=� k��?\za�|��=Z&_�&�Q�/�7��O�����w��V�K?��j]\��:��=�)d�����2.�N�+:��?7��
5ං�t��o�\M�@¾9tt>a�՝�ԤR�$T=\� R���!��!�?"�������,Q�+"�r(���Zz�,�71����
�ڒ)��d��<�ݣDQM���M�R��_m�$�)���?-ݿ�$���e4�;�w1��!):p���J��q�h+\\�ó'�;mC��o�ͮjj9�h�#�D��yO�6�%�V�	�C^�5'M�~������~�"\&{�R@�J����*ӫL���}��a\	��q����i������ɹ��n�k
��;��6��8�ĕ���ևc�n�l&�KQ�J'�O=	�IA|?��~����Q��)�Ł�Y��#��Q�Y���t"Y5���Z���c㶷,�
��iWq�A�uWD&��0��W�T������A��QsJj=��`h��S�m�{xDr[�K���`�{��&������q�*��ீ���C�w71i[�� zh�#���IZԛ�P���n��+=�Bh*Y5�K8ip%�%{��If'���r��y��? <���@k���e�o�SA̼NM}��9�+�Υ{�R�Z鍛�}�@Ϗ�
���1�,�����A�>�M:W̾D5*�[��sQ�/�K�n!mM�n���+�&,Q�W�}@��T� q�{R<�1'^��y�)��w3k�4����|(eAā�:�sC~��:K�	T�[䊏c�CFi*VkZ�?\4�M���C���3@zj�	n�Eھ2����?�T�G��U�-n���=T��H�_�\���VV�yq+uwC?ｹW���`�]"��F��X� g�J�K��@���Nᱵ�> �	޽����#:�|���m�����#���v�n���H'v�L�^C�1\�241]6�vF̚v4�ΐR�~U�8�\܀0d޸8�1ـƊ�Q�6���ssߡN�Uk9��
�����1Ǟ�ŷC`����g��9��PF_c�i�3�C���偮G���-Zf��m4y�HY� N���͝���هHMH���S.�s�c����Z���8�Fù����ʑO��g}����ђ��/���Őۺ^�5#V��˼�Nlw�ivV��Ҥ�"��r��
][[jw����ɐ�%�x��h'�,��@�*�'�lII���u�]��� �FoF���4�s8�!spo��|`<�U�J�%��Ϣ+����
��Խ���>��e�
[�tv�o�ᶈ�e��=%���/���8�0ӵ���/��q�:��EjNB~��l�צּ�y.���J/�3U��i�< �-әj�7a��ԅ9sZ�
SE�f�A�W�~�r�Y	�j�Z?)�N/&��S7�E*H,�ã�wn|�h2!bz\R�?@�+���[nhV�x�ɨ�!G�.O5�̇KM����Q��ܥ�%�e �Ur�Kk�u����3��?셽I��d�$�_V[��s���� �xl~E�Ip��]�nBk���L�˽v����)�u� ���wCJ���ӕ��L����-��+P�%��I+ȕ����Cy��}�L���@��5gV�CA��e��#4�n�[��oe��wj�jbXoLk����	��7�t.9��X6y���ہd�ʃ^�)X�C��.K�C��*j3�Ek����ɍ��o��AoYӈj��$)
�{N�F�Z3Sj)����%�$_F���\�~�%�_%���q�5�w��=Mx�x�u8ǈj
�#�j�$Bo��4��[$ �I����W�*��7$����Ѿ\���X	X ���@}�)3Q�m=�C�t���B�W�Bxzq��1��M�����<����&�:��o�:*;�c68|тy�ez$�AN��GP�C�$E�o�Ԭ)�����߱�������I�[����r�\���x|��,���WN�
�rk3V�͎ݿ�Z����쌒H���U��LN�й��S��q(1�7@T�#�tc�*��ma�|��(����`R��2c��ehD�l���8��>p�����<p~�p���E�D�E8�9�T7.�S�C��	t�	� �莤�y̵8�����&�5U'g1�g�D�.��
�l[ʽ_�x���̄i��m�%
u��paz�9ٍ�G����-��#�C���/t���{�����H�Wo�A�N>���Y!_k�ǫ�	+(=<��_��6�l�g?~�I��{rB��C
��H�����9�r����DT�=I����y�m��x.랮a�v) m�K�ud5��P��#�jWijb?���M��r����)�{�a1��J)i謠O�\����?�P�,�l�n����OP`}3�.�͟���ڌ��ڮ���a����bP���'��,��!,�Nޓ�#�'rm��p�K��Ŧǎ��>��xpk{�O�,5�ε`��h#B}z�.�8��	A�l/1���J�X�~���cW�$��⢵�P�WE�j�0<ww(]E|(\	Wq�k���0Y/{��ӯ�Cb@�$��ޱ�Kh��l�*��8R(��L�x}���ʬ������AA��(��[�
|��K����?CLΜ��d(�!Q/�{�$]'F�$u����[���b˃�6�C�@�kwm��S�I��[�`�Z�=��X�S�Q��%�%ߵ�����_��\5wkZ�N�F�K �S�d��_���@v��z4�:��ouG�E�AU�	���Ʈ�������uzՉ��/F�L�=m��j��p8��M��]�I���V��V��c�GR�R�?��!��Yd�4mGC��epE�jr��ũ�>����.�e����OFdR��潿�ŌC[���0��(c�W$_S�ߋ�p<�gEK\�7���t�K{eaP��_�އ�2�6�Y���v:�%c7����-1�~o�Xh��$Ed��T����Ӗ��v�N?�{�A���t+g�f�3B�� 	�x0��5'1�$]P�F���p��?]qȯ��m��K]�"�h���5�N-j���e�$!����w������@�ͪ:����t:�n��Tq�@�� N�?���K�r�ޙ��Ş�*+�s'����<@�=۷�^HD"G�����Ob��R5>OXYPJ������^a�N\F����!������%j]�f+E�C��Z�����@2�bP֜�@�>�̺�����R��䪮7ײT����"-�G�����*��\��5l=��Vp�H�=aNZ�;e/R�sjg>8��I�%QoĳՆ�Y\��Z$uNc�9��Tb�m�^����*������꧒���<�U_�"_�;tG�W������/�G�@�s�`-�8V�SfL��M<wMF��N�P�ރ�U���^纲[a�ѽ.��*�����)ʆT�����n�P��KAs��N��d������%����k�,+���qB���V�܈����VO%B
|�ǭ�kA�Si�{★���0�q7x� �,�m�_��ܹ��  ����wk0<K%�-�]�~[��N���ΤH�̈ͤ����a�s����n)l�`���1 �}Ԃ�v�ʜ��F%�@k|��*VK���i�l���s��p+����1ō��Tw8q03��v��R�UӏϪ>Cp�����t :w$B��U5����#��\���8�Y�鿝��u�����Y�2^?�ߴ�?P�ExX"|�>��3��yuݻF��M݊���"Uԍ�'��\Jz�?a������_�9Ι]F����S7(������&���(b�p�؄�=�I����R��f;�V��cj����	B�C9�rf�u���|Q<FEw�m�l�!�����3~&��rI	8m�����Z7O�|�^�YX�{����8�g&i�]�G��yyՍ��ɺQʎ~$Pz�T{�`}qG�?���	����f;#�g�4w���(�!ZJ�2W�&����.J��eB�B��&��s�MG,G��gYX�|�����9:ƳS�L���Ʊ(3���'d�CP+���~�,�;�ÇR!��]��<�N*Ǧ��t,�������B��C8��d��v���\턦J��Nuk!@d�7��v"��8F㬋xn���*�9�O�2w7h�vt��7#���I�KzKv%���_E����x�X�T/Va=6J��eh��*W��~�%:]`��=T�aZ�������^}��t��DDz�LYc�֧�T�����+�
��BB��x���u5}�?U�io��mP1�b�m��?K 2���a���P��5ٚ��n:�P�rr,mP��V2��[GFeD���y���I� ��G<�O8R��7�3��+�����M��i<��g��6� ]�D'��I%��+n�� 2� Vw�V�� {���=ԅ/ >�E�����X0�ץ��w���Ý��<d�9����H��r���;���#��|�>@g�/�R�|	��*���j�W�ٟ�|�S^�?��W����Sd|���F�i���@��}
7�0xͼ�fwa,S��g��W%c�1��A�n�J��θ���Wn��x �މ*A�]��@/�z˝1����RJ�	�M�rL�S��N�����Gc��C@n	���x����V%�s���S���Ӽ1_����0lK��jlhEz x�Rd�=�!�b�K�Mpbڋ�S���O�:�2���\�����#�-���#�d�I�����CتC/�`�#ʍ��%[��p[ԉ��%�TX0-V"�W�qL��sl�Va���y9e������CZ��QfDF�j�8���|��a��x.�S���A��B��?ݽ�^Y]�s���Z�a�gk4�czݰ\�l��cP )����/|�p=��1�-�[s��̣�l�i�stF\K[���:eϸ6	X��#�m`�������/��i5���uN��"�U_�Ձ��18U<�E��&2�d���.^��S�ff�=�I�*9X�C�H#�4sB��FDq��_G�r)�z�x�E*H)����
m���>waS��T�$�Nħ��f$�u�Qm�Ⱥ��U}a�	�� �v{LO2tf3 @
�ze)�<s����xi&�D	L�߿[���E S!A
��̜@ޘ�ؾ�{2p,<2��U�����c��]:Y3��r�{��vc�����;3:�z�&�=2u�;M��[�ШE�n@^�9T/�0�8�Q����O��C��Fa0���n��Y��9~o�u�-���c�K��w�*�����T���J�{����M��IM��M+�x�p�'����o��/n���I�||�%˯��0��X�D�c��$���7N҇~E�
o +���[��8��{Ni�/��ъ�'�ijIm6׀d ��>]���!d��Зsd Bؔ	����\-hD�J�VrQ�Yn	;�T��<��tX]�U3�|�>��n���w �|�f�n�3(��^G%�*w��IrA)�0s�G$U���H7�s�bU�l8���x� ���乃5��ц�(scx�>�fn��Y��_K��]@W�1o{ly:e붜�p�-��v&�e��ӿ���<��|��?3�f��� �l%Qn}�W����y$��.�,��tAU��,��/�[b��g�(���V-�G���T��V˯)	��ɦɋ���/���}������d|�֑��ve^]UC�F`L����P�W�1��Ph��$ؔ�{0�� u�`_3�la��H�<�Jp����v`5��<F�"�j��&����fR���.�(�?���1n�!*:2�P:�YX6�tƚ�W���ѡ)��~�62��[����(Zb��2!~*зZU��Ϊr�)��yg
q� �2.�%�=Z_}���Smk-�m��XG���#� �Y�*��2܏Œbh�_���C�b��2aِf�y���/s�ו�=���[���X��VC�w>���J�����]���֠Q�Pms �{F~�PA�Q�:�,�B�ŽXY��s�ж�c��7$(��Z;{3��h+��g[���	�t��$�s�6���[�N���ր�x�;kBI�����D����ק��i��#IL���a�x���1��IbE&���~ ��3pp�A��N�nύҙ��	2)�Vo��-<;�E%Q�_�	��.q���ȝ�I΍yO��J���} 5V�k��Q��L܁2X�ʖe�{Z��3��fPc�cT�Q�6�I�֯�)J�?Em�/8�h�	�Ƃ�E*]&T���0����á��Z˿L�����%�O��e�S�!�	��XQ%!A%&I���*뭀/i��KX�>��(���_�E�Iœ�eZ��i�_�D8�N�$�Vj�]�_]��3s�`3fW�����E�21�:���1�~eåNT�,Z(�(�hp��}�����!ݩ�!�8�̉d�%��%Q7k�m`�ms;�Ҋ2[�x`�0���X�^�+����Ӹ����Zϋ��	?2�,�vcw�>��R�2/'����_Z���fw*}W�R�5|EYu,t1��A�2ku���w��G:�v~� 2�~��)Q����s�t���l�ZS%�'<4�+���c�M���o=ù'+@��Y�I���Y��8hO�1� m� ��G�IC�+	��K$=*_(vd�fE��u�t��-ob��ړ��D�����|?�ߑ||X���k��A>���:F2ccxmz\�~Q;��MOh;3Az^�4�q:�D&�x��:�G5�L�m�}����y��c\��|���� ��T:꿨��4'��,��\��!�'�p�IJ䅋��e�Ԇp��;�0LV���ar.������Bs:���*��?��զ0����E/�	�nCY2�,6���-%z�|�������Ǎ����+��#��4[��C���f�w3���f/�*(��]�[�UE�TtL<fV�/^��cw��c�f�����1"���N��iulO�)�%8�����1;l63V-�|[�d�l�l9��ɮ��3b��{X��y6CY1�Yi���~�37�����8[VM�3q?��^�j�C$����}�XE�c(%v�{���~4�w�(�9��6��ڑ%�\��3{z@M^y��b�}K��+G�8y16� I�&�D�Jz�I�;U�&yQ(�-�/G�;OF�IsQ08�ShW���qz(���MFaM�%����D?WM`�.��!`�I���K:`�H`����w�9H�U��8�g
r| S�Su,lLQi׶M�'�9���H@ǸFZ��` �"}��9�I�C���������2�̿х��I��>Cf�@���_x����2�)��%d���G�]�$��c���+?�F�)f�$I4���:�6xl�����P��a��^�/qg��򐶯`��@��W 8Аe�k��Vc�c$`�%�����C�N��^��ܨ榻+7�BBl�J����jp�W�B@�D[`� n�@�3p�����:%84ʙ��&�����!�B��&ؠ×�"}g���{kC_� n�(��vʆ�er�}Ӯ� Q~.�	[��wv���G���T��A�°#�݉ >F� �X��v����pb
{X'<���<�P;T/��j����3�^��B�<���}d[OAaj�����:�#�M��k�