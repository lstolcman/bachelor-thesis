��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�0b�:.}$��;��q�y�P	���=�����T�==��Q�#Y��9��? �vH�(;��sg����uyQ� ��	"f(nvd�n!t��A���w�臒�������y��qk5�~�#
(��X�:d�Z{�O�b��*�w�e��o�3tQ�DP����V�Rbx���ޝG9�C�gAb<���+5�aYC
��:�[쨗�H�ĸ��;S�#�fI`+���Ą����՟�Q	xKA�I��l�^�o�%�Jz��n���g�[PN5�qc�M����(0����e.�==�����=Z^3�U!��m-�w`v
�{0�?։����[�_DH7���e�rȮ��O�	�t��mkD����f������S�6T.3x��G)�Zԛ�@�-SK�D�`�kp��ËJ����yP�x^�ϡ���Jr~kz����{M� Fx36��8)���*#0���+�u}x���2��
��7q��s��ҚjJEN�<��b}3yFTo(��1qW���K�ě�v�0�Χ0�寚G2g�:�"_���P�Y��i�
7�S.(C`z��(]ٔ��9�.�쫇Ga/j�9��5�|UQ������vm'ܨ��)6vD�G;��1��r*��[�7�Yg("��PF[�1�F��o���͠�W�����]*��H��v�LG���pk\�/�N��uls��j�H�G�J7cogz�2^:�u8��ط��VP�[	t��H)�ޚya���7|O�P�]|��~�L��V|{r::��)�i�7��wXL3-Q��"����o=��/�8ְ	�!5�@�r�˷���S�<h�dM�?Q��|ƪܲ����u�`�!�
w��T��	��ʂ�f��G����}�¾�;w�|-��Sq�#�LcZhr,�2��q߿6�9�<�M|�_�&��j�\�S������vų�<SK���M����sT�Nh�#�Ks�ȳ�ڕ�b��;6#�3�v�T�wT>�X��-
AV�M�p�����5�L���ߕY_B���<<k6�c�ܜ�n�+G���0Z��������`�c���W$�N��ϫzn}qe:�Wk��\G��]�Y4��
�z�Lw��lB���\DJ/�OK��Mq�hD<i�	�m�#��W���uR!����3	�J�-2�# Y���=������v��颻+�uZ"��#|�X����Z����'7�K:�Emq~�+˵��+g�`Ɯ=�1�c�>��4X+��9��V���!�6Qd=T@"��+T��2���"O��Kn��'��^�fQ�jnI���m�ͬ
��W�y����A�[g��9����ѿ���3��&�/Ml��s$=a8W������֐��y"�z)����t�&;E��<�ނ�h�Vy�M�$2 KƳ����è�1��q��M��k.Ȯ��6uc�>-и�h* z��6�@�.�Ta� ����4��f���==��!��^���t��h�Y���x!�k���v!�s!��8����xz�#��3���pի�M�?B�yS������6-jNX��I���"˝��;|�v .��?hT�yOD�v��[ٮ
	�niM�3����C��`o-���C��a;�@��{�ˁ��2��z�,K%�E˻��J·^9�1@ߍH����*��-G9B)�����@����@��B�F�> cEf�J���U��F>�m&&�]��}N�.P��i���^��W���wa4f|:�W�.,$�y��-���F��`�(H��=x��"�A��) ���;%���ə�yC��[��L���乻)��|�q���ƻ���{�x֬>g��!�m���/����cZDp��4����.�+1�+ ����Z�߱6<
bv��\	�WC�V�v��B]e�qϭʿ��1qo#)`im���S��m�.<c���e��G2���cc�)?{�"-_?Lٮ��|ۋ�E������`�6�V�ũ�����T��V-)Uu�Q�Vؽi!�)�������P�"�ݣLІ�M���°?�O!N:�E���ʈ�H�m�q�,'.5q���i�#|#�"��4r����KV�Wg�z�d�`|{��Zݵ�Z�m,S[7�M��%���O�(ktD�'�T�S��]ȃ�-��MN��]m�Y��em<��DC��IyJyS����z�5���2�	b&u�I�F%�RI0���\DՑ�MY�s]Q�<0Y}�:��7!�7�ob`+5��f�m�K�|���-|�C>�bЃg ���tt��8��n�^Du>&��~��.�^�JpďXd��
�[b�L-W���]U<C��g�f3*>�y³���0�B�*XO�9�u��
@��$n>�Z�!B&rB�(DP�}�k�^O�����S�JΑ�P�����A�N��z��s��y��di�[�'���S)��*��f�[��s1F����D�Mi�u����aI��y��#��3����{��姠��9�pn"9X.�Z���-����~���ڔV�̕c̯��y���xm��ʋ���"U0
���u0���j��5�h���O�!
�Za�xP�laI@��B���pǂݢe�sX^���0An	�\����c�tST��ޱJTrG�ƿ'��? ��ՃWtd�i;�ݖ�|���6���3���NO�0�	E��JSf�9�N>6C򱊶��Cw?^�mkT�Hwٻ"��2AGށ[xӉ��=d[���r�%|O�+/��&54��� K7Ԥ�:��;�l��ƨ�MhSj���e�tFI4���b�/� ���!	��z�f��~�>���kB�Y�̵�m�!�3�<DlYXyw(�WM�o;�b����Zt3k��πl���I�*��Ѿ�O��&�A�0��EF�<�]�5�X��D���ĉg��)x��=g졂ײ�xJ�Bj�J<�8K�Ï�)����uB���o	�1M�t���G��I��8�#9�hd�p���6��HI�N!�·���?��Mg��s�\�M��'@2IqG��-3|�(�5�|HqB$]w��^r)GKD;����3)�ח:b4+�����vk�(��Aj+'s	��x���*� �����)d�F�'n�*`r[�R/t�g�;,�����/MZ�:6�� ���G�}b����m F�F�\Ä�/޹�X�=���A"���_���5�z�#��C�c'�#��#�D���{�$�H�t�9��M��:�Hf�l'z�Fq�Їw?a�A`����F.�����}.`۪�nLf'��y0��Yd���ɀ��zX�h��w�;�%��ũ+�&j�T�G�*Y_nI�Ʉ����¯�K��}g(�T�73X?���7�/��	_��Z���\�q�G7|&uQ���td�eG�"#ȆU�S���a���9�齅��6뭃�ۉ�	�M��'An�*�]�T%��N�'�E����"	��0y�<y#bI���}jAX��"��&r��6�ľ/	�݇����,������ �xDU�td� J9���i�|��5
��F@�h �5��z�|u)7��{�FX�^�އ�Z��pr�du�^�&L�64:r1|R����aL�!~r���&d訞B��L!Zڦ�+n���a^`��QM˃Z�i��|���R0���܍�F;8H�Z�#��m�P��3(=�_ Z�x�ڤ���EN��e��U��W�J>iAA��s ��uAh�;QR����lJ��ެ���OH&���Ltz��)��f�a���>^����m�>*��	@�ߕ��(����F�N��d�m�	��NH�1��Y�J�~�ҧ�Ja�V�ǲu$A��BL�?��c�c-�HO{$ls�ܓ����Cu�dc�l��s��Ν�����e襱���WJ�������f�眿m�	��	.�
�z(�d���k�s����Ղ���T5�HBG �K4�M�N����W���3����H気��%�V�;N�9#f<<,t�9A�]yw��_�ϱ�8�[��� �ڐӔ���O/�1�v��K��u���iZw3�ʣ��e?*%fI��xN*H~Q<g�@����
�e^�O'(�����M�V��C���o�V��1�d�t��̡�~���2$�"R^Ks�G�Nӟn5����� 
2f3.g�痤A�(��}s4��h'���8ggDb���|��	R�;*��{�b-������K
�0�~�ՙ 민#D�P@ل��hT�g�T���^����+,�Q�'��Y�0"Go��L ��x���;��Oq~����>K��ek�<�3�[���"�j��ӌ�>y�A��FsͪZh�@�1s�<ѿ��vt�+�;�Z%_�V�jӨ�c=`T�F�����Xf�@L�@��5�#-Y-����t��s��h�M�,X~ɔu����{�7�X������fr�:1�t�Uds{9���;��S���p3Qu��#�'K+"ل�p�Q��t��b��e�]
djt���3|�a�E�5�*��d럔�f�)��<>�8���EH���0{v�;����evW�j.q�"1���&���~i/������	`���֭�~�wR�� ��B	A�����Z�^7����ʸ�NX�gڞ�i��Yf ?�!�$�n�8*������N$���6��$>}��#���i#�j'a�pX��لib
k�p�PN���@+b����rg~�u��8�H��SI6p�w*��v'mT�;�Ҿ��AwVq��*�ĨI�J���5ٞ�|�aSό\�W{�g�b��1�+g��t]��br5�8\Rn��Ly
h]��)�+h�MM���б��d�i�vF_�E)?��sl6�`��t����eny;��7 >G�@�zѻ�f��In=��pLؕ��
�Ͱ��cgU|��B'��`t7�+���]���E}oA�xs�*ķ3Cɤ�Nn9��]!q��4�C�W
Q�c�z���;B+�s4�2�1���x�F���W:���%�?u��J/Y�ٜ��sT��3�v/`;	�%Z�T$�[ץ�� ޚ��3Q,B�oj@���xV?�~P���F�!�?�Cmn�#@ߊ�/G'j8����I�4�#�aw!p�[��жҩ��&K��~x%���bD�hꘄ�'���Zus!=��S��@�j��k���N!�=9�fZ� )���:�(]�ux^��?C�zo�>$��������r({���k��
�tA;�f���&�����1x��t�̥��Ai���G�ی��,�#���s����$��L�WPh�ARϧY�Ę�Kx�W��%O���<�Nh*���=g"b⑖���a�'���5	�߼���	'(�����s~�qI�K��S#���[��Pb�;KK���ɩ;�ab��'��A�}ԒK]� %�3+@��C2*hK�N5b�̎��%P�=ƅ�f��B�#�)�b�c ��P�K��%v�pN	��;U�@p�K�/�����:?�<T짌~���@�g�T�`�� .�ƃ� 2>�z`3��'�� ]_��}�>��Ȭu#�n���|_m0?&Ȥ;��wʴ���*�}ʊ���'�?�����r�"*#����z��4��\�&��o��G�� �-��
z��HqFD�=0��~�pb�:@�Y���JXvE��6/����]�X.��/���� ���Q��:}5�?��C���R�a:�ɗ�m����o��/v�A�,㌗������tM�
�� �P"�ē����G�墊���F�Z��$i)�ɜ���q��_\�=���?B
yI�e�m�[���R�m ^��<6�rF���f������?��g_��B��fQ �P:9��`U0g��Ap!]8�}��ma��ඈ� �&y9�n�=����=1-��}���o�4�z�V|z]��TI��#ZA���L/��T��r���!d��N+1�(h��'�C-��Oc�lkkn
<)�ު�1 ��UJ��[!$�ϋ�u����"�yhEZ�J��8�T����Eh�����ͤ�H�Oi�F�XF4����M���(�Q~+=��%��Yd�s[�$:�~�3���v#쁡�����}��?�.�,�̏���QC����_t�IE��n��ö+���H��?G�G2u�	2��5qL����A�k����
��S�Z��u���U�#�d��h�3|���8Cê��a�ľ�˟�Z#�"�옐kek�rz�C`�pϛ��q{��D��1p��d���F�*��o�4ev�+"&Ɋ�ِ���-?�Ts�}K�i� ��$g�sn+��k����N��!!�/�V_���Ѝ?F������f���gz�#�mz�s�ThQ�g;"r�9��V�I�2+�qJ���\'���*�����Ç�����OU�s�-�O��OL��쾷V��� ᆳ���
T<鯫U�I;+x>�R?8QR~p.�r'��9Ǚ�˴�� Wu��h��O�-{H�.%f���6n�׊��*�ܤ�q;�YY]�Z�`��#m���.#�c�[�ݙ3i��[�O#¯a/�!3��N�=���x���i!�ą�#T������N�����~�kq��rC���#r������C{
��z��į�	)kFwy����u�۪�}���^z1�ʜ&c^f�䀘��Aܿ��!4��r��H�~��K�-�\�W���/�6��M!/�b��'�:�	�M���}���5�\7�/6�W�+�5��k����/��}��V����
���P�RA�ϫG��H���P���;�;���bu�6�9��r��v&�� vM�!���z���ZC[��xF��o������b.����K���$���AR�V�u5$!�������
N7´&R����"ʯ�>?�ͳ�߹(!�%o�A���2
�Q%#���%;f���^- b3�190߼��A�(&�Uc M����*�)�RؖЀ\���jTC�BS���ڀ�/�М�vj�đd9#$Ug7Oh���߉�t�H�}��r.i��y��rds4t8�����P>D�-(m�=�*וe�������4dy�����r���?�r���L��7VD�d���i���z��;ی�1��i�B�<���b1��
��+��aנٯ,��ad��4V�@�]�o(�rE�Æ��/�r�����}�L�G[4�����h0���w��f�D��>OQ�O��3�&k�`~񲑿t�;��;� 
�V��Pۡ�c�!��� �9�oq�y�8�Ep�g�v�@���6�Z����ߛQ���u��J���}����pā��*��3[�}F�/(#z��~��hd*[Wʟ�c�I�����O��6��7Lw�Z���Ĵs!�1��E����ꉎ!`�ê/��'�u�~X*�B׬����x��K�3D��u����ݽl��緲��Ҋ�J���ǿ}:���!Jb�Ǽ�9�s�v3��TH!�$Bi�[��Z�~͚��#�:�B��hFZ@�E�C��Za����'4�,�� O_(�j��*	RT�9R,�9\�nz,>�I�j�i�Qg�^1�eGղdh����5��<�Du3�}���m�����l'A���Ҡ2=�f%O,Of���`g8g�unm�?N��N�ץSøa$s��p�\'8FU������c�:�[I�'#��FC��y�n�)PN�M\��+��{�m�|�z�����b�&LJ���Y1pw�u�����h,��̩����I�����?�\=��n���\�EQ��I��]�umW!��-�bN���.��ϵm�!�醒x�^hш�텔��RC�Ĉ�;���#lSQa?�}�e�z�R�\�L>�]: