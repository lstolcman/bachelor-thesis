��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J�-�4ϼA�xu*��6P��i���?���3�Rx�Ct���Ơť��dKkAW��.u�����"Ѱ���8���y~�c���o-=�S(��Eӟ�uC��X��IKb4c�,�C��N��h e���j�giC�R@ 3ˀ�un!�>��<���;d�aj��&}S���j�0.����F�hY�T�c]qGGǡ{{�H��]|�WEW��"����Ot*�p7�&Ю���i��z��Ń���>�-*���I~���%�5�ԛ�!>\�)�a�{K�� (rӵ�}������:��aXџ�ŏi2W��Ss֐[I�,�fv��\�h�eu��x��R�A�9���d�ȭ��k��5� u�֔ Tf�۪���,�A�z�8�z�8@#o�E�2e��ȟ�օ07����9PZR���ޯ9~b��M
��(U汒5��w��!ʑ�Ad�( QA��`۶���_%�#/�q2�j�����3�B�N�ľ^���|3J9Q�-�S��2L����tM�֓��V��cf[|���ٗ]G�����u10z$wP�����sj��Sg�d�"�:E��-�/<�������d�k�����<��vއ��$��V����4�T[XϐjE^}&W)q	����r��	�?��i�:�d�����������`�\������Tz���rR�o���]yu6�����sG�Az;'���v�����d�����A��<���Ӥ;�n"�҈���Ck\��׏~l��X���;f��$����&�����4�Ie�;T[GI(n۞����Cs��y5�-cF���L� �_��T�g�6��X԰b������ ?�Ͽ$D��J���T\�' |����ca�Ooc�%ׯ�G��d�%$���HnG�_��^=�������������^ ��?IB�G�eE��t�#X���n~X���x�w��ڹ����E�e���>�<����Br���GⳞ)��,E�/۴��h����:�h>4���� |"�k���V��`r`= �\:.h
ǪHk�}+u�1��5�cW[�heD����,����DӏŸ���I�S�g[�����B�]��0>��-Xa����?��9���4)K�Z9/�уŒ�k��w��{��h�������qt*������������8��^������~)�E����U�[pO�� ��)��v�#��}���=bM�Usk�g@$=I7�@�1���b�_���^g�(0���-[�4N�^nw��NI1u%�tGhz��S�b�/tH8�|���U��jC�ƪٍ���U*u1� �IV���z�����#'�#�E�W�	Zd���NkZ'N{�}Mƫ�t�f�i��{9�s��;�P_%�������ȗ8p��{��t@Mɽi���y�k��p��]�^ZD�b0���Nr9��ݎ��d/3dw��L�ǿ �]�P0՘<���;w�����^*ȥ%sg���=�x��~6աx�$C'2s�.68�����g��K���X�P�4�����[_�\)��)��{ێ$}��~w�FN�!���mU�9�cq&��l�=��Ҳ �0��TC��/��D��c�g�]��G������)U(��-�?i�=.Z�6j���{��2�U��R���ڭ�^;� S��<�r��3w�h�|���5F�����P:�xD[zSe�j����(+��X�8OC�3�� ���+Hx%���)od�Q�����׌��?��ZM�m~_�i7�E�$P��V�-pt��﷋/���Fr�����bC��Q&�Y}�Ӯ����-ג�}k�ؘ���ˮw�X�C-�S��8�2ͪ������t��/���Ue���(�,J��ӔV����K1�hܗ��Eq��2����o��h���,1�S�GL�v.��贶�h������$ku|��#>�b�RAY�&������^
��`���Q�0-#֨�m�	��|�.��L�o���n���Y��ܗ�\�tY�o�fܖ
��o�:�>��T�����[�w�q��'���a���,t%F�WClG�\u��ܮ)N�">��N���$�ά�s��w����k!d먥����%��ב$������������������L28��7��
�����l9Ld5n�Il|U�)��7d9���y�g�Så,_u��[��C܅@\�����e٧���IC9�/�T��&�m�Ԯ��"gz)�R^�=	J���G��kO�ࡂݑD͟a5��뿐D�?W��O�/S�N�`�w��{�J �\(�G�U�ڳqW_��<���F}�l��j�C�H)ޞU�[.�I:"����=����˶0�faWr���)����S�3fQ̀�+˓I,��P��R�������Ӎ��S`@ǒė�_�"����jo�R����-юp��Br��n/>g$��׹?<�ZT�9��H0��\b��Yy������&?b�p�ắ�a~E���r�m�-����dX8Ԩ��3�u�l���&I� ���K�&��1�̉�t�Wo�X��~�����n6q���̯{�!k j��fVV�[�fb+j~����g�>r��q����K?CN���?���\Ʊ�i�}Ɵ�Z�/^���甲uX��P[�����- �z���9��� ���p%����u��>�ӛ]�C�f����*ȭ��D�K�`�L�o�B�����)�oBt3���#���.��K��%�%�Q�~��S�T{���*�0�H~4ջD`�9��3��ߍcQ��g��0��J�c��0!�G]�ѣ��N���U