��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�O�5t�"��شV�x/Tj�T�.Vw�3��oO�����Y�4�J�E����8n)t@�;�]붾DJp�cG���:����m>�(�P�+�4�r�m=<Gү��T]2���ɚڡS�`��IX��I�����{-��LOL�)���	��to.��	*�8̭�ȑ���0!f3k��#7�phY�ß�<h��ghW{6�Ira��p*򐍕5Z+}R���b+1���a<��[-� �!����l��`#����U�f���;���ڬ�0��|�R���7N	L��'y�����щ��>T/�B^v4 �-鑜�
��U��x�f�;٬":`��Uy|�W���Zў�n:s7_Y�s��/N��?7/U �dk-�t�a�
�I�tY8t���*,��$�
i�=R�q�hϸ��SP�h����
�x̗��y����b��ѻ^1��k9v��n�~���ގr���f�;G����r=��f�g�n����O������(_'hڲ�2��&Y�2��Q�w#e���_<�gtJ�p��´B<�y޵�Ie��Ě��i����K�������� �FjU�ۏM�AD��XB�q��e>h�mi��Aw�#e�`���ɪ
ǏN�V��dU�+Kc�Lq�/��TuM�<��Zo���y����ď��4�����B���z��{9��n%C�:�fM���� yP�!��6ڒ���
�"	V�k�����WS����-Bh�9-޽�x5��xH�a!�}dY�+@��vc��i/G�Go������?�!�d_���܊�u���w�]����J��/���L�W�3)e��X��1�O��wSB�u�"�!;d��D<���"yF�ig�zgPW�E�[��S±\W˾HJ#CY�}��/��0oQa{�;��;C��v�qX�h���ɦ���֣��*6pv�<<0�v,�_x?6x@0Y��=�����L8R�8s���O�D�V; &�+a((L��C��� ������K�>����������XѾE�'x/�B>
h�:����E���2�i �/6肩�1_a��{�-�=>g��`�{���l�i�&N�V��H�M��YJ(	zi^#x�"u�I̔/�w�ԙQ��C����}���&�^�)��M���f���	�oji�UX�I[{�5=؅_щ��I���$��������p�Uk�о(*Kd��m�P�v{����cy@9#��ږ��O.D�a�����447iڵ+LH�,�.��G�-x�x�ޓ�lס������I��s��|:.��|MR��@�=
��^F사�\!��fkhR?���ouRG�1��^C�
pk�I�JMv�p�ŷ}�O��n�4�����>�)�S�_�f�؉�.����0x���j#kAe�G�mV��g��\ ���v�x,���~��� �ß�跘°�|�������tV����e��9}7�jK|����0��zGV�:�j�
��񋅯�����Ч�(k���o�g������""F��1�R �D���hF0���L��ڳT���-8o��@"w
Ĵ#�<a�^f��+0�*���l�9w�e�6٭�l��2{�&���y֛�o�*_�bt��%*̕�fA#�:�m�97��e���(�6|���y��,WN �o��YRΐŹ��Qۆj�_�)�]\��[�b�2��V���v�Mt��8G�6�%�(U!���XۼU�q����O��g���K�9�7��?�܁,�<�7��s�8�����`i���Ͽ+�h�(��T�o��3���,Qݠˋ�w;��"?��̶�=ˁ�7�E�d�U߭���-�3W��Q�x�u��Br��3���gک��K�����^�P�
تM�呆z?��#^g��/P7؃N��1��?����n��x��MA%1�N������#8�ӐN��Û�%5�M,��^�7�i���V��@N��k?��(Th7 ��g&�]���c�<��脆-�oV.0Ӂ,�,�ORK_���`�I��)��u#���D:�S!ڸ��5����]����<aX^�G!�]�~=O3�B�*$#A����,
�Zf��l���D�nE�\ZVy:���i����5�%2���}��7�F8'�Je,�rZw>"o�7�f���������^H�}]�>0JӬqr�����B\	�#G'��W�Y���4\Ca+�wf]Z���1�D1J�4u5�������X�u@Ԩ����!E;zdl<�v�T�[��2�"^)v~ɺ��NY-�CpU������T��|�Nirè��*
��y��[O��vj5g�)�� }��|k�T���-V��f5s�u��Ɗ��A
'=�£��#"�OF9�K�ch�;a�A[G  '�9ޘ���&��=�c�!���2�F�J�G������o��<��{�
Ѓ��Ejɚ��8+�����C~�����e�)PY�,�?���\K�o�M�眨����'�x�����W[�M8fA��h;1W���%ʶZy5�ZZ��#>�|�E29=�,�]�d��օs����� ���Zz��(�yc˟��Ff;/*Y��I8�6!j����}���9ڳ�І8��"";!M����Z�)����{��~�F誴?�4�h�;�O��@.�mBA/�
Ѧ�e��&�(Cx�. ٷ!�����B}�~K�H��N:&�yh2�kf���ɧ�	��90��=��U��U@^����__m�B��$��8�����H�cӜ�kZ�mz�Q��R�^/6�o�4æރ�C4�O��N9*��F��Y��_���d�e����+��ƏX-i{���+䌒� ��~�6�)�ԙV�I���:��#te໲g2�Ķ��B���G@KF�X�u�(�~^{<]vc�u�Ze{�i� z �}�m{����Ϥ~R��}L2���ep�
�[���)y�f�X���3�%&]E@Uۥ ��y��]qfEݿ�H�b�10d���"�.i�eb�������]CY�#p�16�[$K1�r9ʢ��c���2��4��Pz��D0���yvP�2DM��8��4�*�E�Q�Ff���J�Y:f	W���)��e*��~S��62u=N��A�7l}	=��U/Z�ޫV�`R�]�W/�"��(�(g���=���my� ��d�*y���^!�~�KF�;�`��\�H��^�0MV�*-�#�Aڢ*%���$�Q�@,1���X禌y�P�U�u<�8q?�9uѬ�r^����$�>�	i��^1�*䨘��0�'�~�ퟩ-a�Q���4X��੃��o�ĿV�phvP��K0��ly*<�«���C��r���(��*��Q%���
�@�v�3���Rx0*Z(�e)׉��A����v�Y\d���뉆ύ� anK##����e:~w���b+�35���EQ��X���h:LFc��cj��[h�/ެ*�ؕCf�T�N@�QM�j:�8����^���5�T�`U�m�x\��1��#a?6�Y�O}�]�R����_���P�D�߶_����X���� z��;��	s~I}oX����\O("_����r3T���E�X��>���~G��Z��2�Qf�}q��d� ������sAo�	VıqqL�s�iW�o��Z}ipLbr����Pw'��	Y��s'}�yn�&ͨ�Es�0M�=$��Eޠ�cU���#����Ԍ�]�-�0�I�|b�m�!�:�
:B$f�mŹ�
4��,U���f�"�[]]����t6^�,殂��Ÿr�������d�yk.F�}����\k��5d�CF"��i��h3����6���&�H��v?J�j �F�}�D-n���ڪ;O�ԭ=2��}�Kf�tH��B��dN὆ �˫����H�%�n|Z3��qc���n�B_�0a�Y�̴�| ��O�QlM��(���B�A��U�9&u��t����4�� H�(�Li��5OF�X�K�~1"��H��4�5~�Uiv*����B��6�R$�OO*��?�߈5c�H~U����3Z�a�!�0��cX(�t+�MC�o�O�G�����#w��9�y��'��_�^>�F	+9!�
R�c[���R�69?����4��@�#������OqN7-UK�+����q��-���DO��G�=Cg��Ԩj�~�Xx��64���/�ߕ�����XC9\��q�?1.��2``�D�t/��+�iH��Z��a��e�$�"��U���������74�Br�ϲ�OjG�ۇ9�B��ile�0]��W}r�Ӑ�Hf��C�oTN�i�l+���jOKG<��c 8�&���p�N$����u-z?�t�Ii�L��Hr)�V�өx%�fR���o���>�D�7�#�8(�!d�k��uG8 ��	z�0g(�p���}J���gU��Φ�\�>F.�}d�����=9o:)�Qz`Ŷs����V�DɌ^��3��:.-X���K��wղrUt)�Z�(�ZZ��F��6wnLȚ16y(��9[H�k�zõ�N���^�Yi2/��,R�s�8�:u��9$\�����Z�7�F �(�c��o75�=p݆lg=�J ���4	COO�4Lrr�+Y��P�����F�LPW'9Ǵ�H*ơ�W��o{ir�b���&�[R���/Y�7b�==g���]�Nw�^q��z�ZK��(BO��B��P ����.���Cie�q�\�\�&���ƀ�;���cҴ���IajCω���~sK�Zj2��K�ռ�B;��é���r a����tT�,�!v͚0G1b�E�L<;��$�K��	hs5C�51��3J���Q��Q�+�D����ʻ9<���7u�
Z.�/�%��}�[s�3�)Uv#�H����2e:��y�
�Dl~�y�=�s��a����v�W�bXzS1��B�sRع��PՇ_���5�Ί׶=�-g;����S=��Y���F�K1��i�'3c3}���� �� �'</T�s�K��F�WΊ�vc���j�� �iD�t^^e9Yݨ��r����jCme7v��͒)�h��IF�{�P�{��\�����dǑj"s;K���B�z��%m���ʂY�{��9��WU=��56D2ԗ|�_���Kݦn~�do����Jf�|%A��)��~���eړo�V]�.�L�݄KF�S���'<tg��
�t,؁Rsy�A�����dP/���=�t�7}�ʀ��װ�����ڠ��	|�Y�{���YԬ���d.}�#n�4�:����{H�,[�\f�;��k����M��C�\sPh`*�`��wh8��t��vu/rȘ[������9&�o�@���J�u��]:0A�>Ǆy�ǋJh�LrP:�1N݉�!������u�o|�'8 �D��υ�B/qt���lΠP�@�&�����CV��ʒ���zݱ�A�Q��<�F���c�}�L�o�NE�!����M�7����GKI=����5һZ�c��p>m������jxE�!E��b��B$=H�j�F�\�� �F�5A,t��*T�:���A���Un��ga����4�s���Ћ@CR`"�d�Y��I���v`i�DQ��� k��.�j���~@�����u���}���`������4 VO���ǒ�N �Ų�����dK.0ACʥ�� Lĉl�p�?+�B�Q���}8�P;�	?���RV>ʜO<~'""nIy��|�1`F�\-3rnn��ß�]}8Iu@$R4�����%-��,Ac�lV�|��,�j����jĂ�o?��u?���J�^h��E�s�4mF�K1�k�
>L�������x7�2��=�x��ծ��d$�|�3n����+���W����+V2��47�#v��x֖WQ���3;��J����՛3<��Ĺ�9sb�ۃ�������]����Y�
���Ԉ�m]d�y$P�?4�qI�[�}#*��<��:��/�C��Ԫ+!ԓTɻ�x�6�q!V�1�4�Δ��3�حY�Rr?�#c�_�`UQ�D�`ҫl�'�橡��mQ��:B��͐uަ�銣��x�p�!�¦(2pt/���	e�T`�MU
�I��'1�]�C~���Zg�c��	�(] �,���@l�'�B��f��}�����*�[�M�8�����	�Z��6�M�d�]�RY���XY=b�^�τIP�;A�濖8��l��,�boW��b���ʸ�����V��JH��G��:�M��%��?&6�}�Õ9���޽��5fl���:\��[e������Ś�O���k<����16�Ͻ�SE�.�;�l���rKȋ��ޝrr�i�ź$�r�]̘uq�֩�9��M4��$
�){g�v��i���L@�4Β�}�j:�?U��N���#?���g�QJϚ�1ZyϪ������ʼeIf���g_��=/to�/+W{��P�#��s6�:�=܏c����f�n��C�H�0l�&GN@��@5�T�B��!h�lF�^��*���CI�}L��H��H |�[$����WI��t��?�c}ţ����B� �x������.�}��Δ����_�D-���F3\�5`s��޺�N�W��}�lÐ�{s��잀9�H�?n9�wT2�z����qBYC

\ra��Gcw�i�90}��Y�¸��������Ʈz��[��g�b'�U|>�#c�̌�ˡ�"M�v6�=��F��T����~1\ZX�pqQ��M2������mc���{+nS��j���lJ4�����s7@ڰ���Q��z�}Hv�<9���^.�]2U$��!���q�O���KU���^��.L�����
�O�+�~����iY�S`%�p��֞�b���j��ݸk�.0B���tx��ù̥�d� 7'�~�А��EM�r�Φ����Ӿ>��/�(?O�D�G�Sd�?d����2��L������؊`���F7��g,aXçCOb˴�k27��	%�P�0��a��T�o\��h Z"mC���J�+����L��
�J���3"�r�ȍ���Wc���27������i��VV��9�#I( �k�6�V�z�yc��g��������"�q���͍�5�.���ލ
�~��z�I�,w.Z�@l���5�r�`K�ANA�i� �5.jkg���_�$rR��I����΃�iȧ��q�HO�R@^���qX. �� �]6f�(��5��G�c��	��|��.��5���^��+���2�`��n����cH�ً�u�m4[������r,C��-:dN5W�ڪ-|Ǎ�L*��>�:�ǚ����Ofl/�(���nVx�%v��m��'�!��n?x�X ����-������	*��I� F�;π�2ߺ
�CW}j��E!c+R��A�P����wy����#�� �[��.����NE�LZ�Աf�����`.��1�� ��j�f�i��|�����~E5�Ձ�|�ms�x0�� nɬ8�#Di��E�TY6���d-�
5��'^���ҕǈq
�3Ȓ|gZ��(�*�?����Gz��FU�7[)M�����x��f����y��.�Ʉ��-N"��(��[@��p /<�!�!�F]�ڂ�C������(��5���r-	h��E&���q��f��/� ��}��w�v׸�q�bgE��x'�/����Q0��
&���i��*κ�v��x$��4��ت����h:�hq'���o�5�)�a�0����Q3��#���lK�p(��TJ"���8�H��&2�������iǭ����ZeΈj@�,�jv�	������c ����~l�}�s]
��������sg�?5�IgcN�?��RWm�!7%�[Dw�.�ao��B�	T�2㶽dM� ��
���o�O������0k�|/����
R~<��ɻ)�h^5�j���wpDTf>W*����C��\�K֫��{�bACO��3��q�m�j��_� ��ۦ�/-�ĳ
�B���J�ZSv���&	����hLQSo��0M�.
���-�G �_ Y��Xʪ/:c�?v'�o��
�lbo���ޣ��
c b<h)"��3��.:�ۃ�k�9�\R��r0RT}}�$��\�5K�2S��_V��#�1u��F����b���qQ����~eM�>U��s��6��[��Vm��|ɤPqﴅ�ۖ�=�;&��{8���@B�<[�I����V�M�+�.��t@IB��G~ ����~��/�>�ģ�mXd|��;�N]�Y��|��%f��X����Z!����"m�y	74��$��)���������伻�t}cV�;� ��Y���a����b�.�ˋ)�
�h�έ��r"����kon�<1��bޑ��@�P�h>�m�x�d�T��ufp�`�܇U9l;��b��桪�O���Q�{J�5>����[ʀ�V�W	�h�m��OWp9��Wyn�no+(.��ŷ��e̠R1�a�x�Z%�"���A.��k�{
C�I��X"��F�Q�8�X�� ��C�X�q�nS�NC���{�A1PW�^`����xu	�s�#�<	
��0��w��d�J�G�a|J�>Ec��w��^Z.|!��M�s�37P�}�Ӎ��&^��3��8����گ����V3��i�8����C�]�}$�tm���#6J����a��g5	_�����~�H)>'p�����v�=u�pT���7j�^�"�h���H#�S�b��U�B�n��-�n��,v���p~����m���)V2C���������a�W��z4F� w��􅂣�ǩ�Ey:����0^�dq4X�ao�k��ߚ�6_/*����gPG�\ E�ư��r`�#^J*��hx�?�M�W��d��:p�7~��):�;�J$�o�x��F������i7�t�k=�	�u���O^�����qM�9hw�-И88��#����r[�i�����:+NۢT�����*�۞1�@�*�X����Y"]-#����N]p�%}�QK#�;�A�NOH*��@siҢc�/�G_m���7ť��jN���I!�|�1�G��&h��ь�uX����,+��az���bOb�@0o��bs9ÍtS���t�E['x�P�g��9'.���"Ҍ*|�KV��+�f�P'�g�_ˑ-]�Eԍ�3��	94g�m"�uD��k@��zM��]ۯ�;�k��'k[�G[6�FvNϴ]f���4~]�N��X�>U<���J�h�2�m�2 �$k����X�w�1���\���;hP�� xvW,$ߪ BAQ�qh1(|��s�ѯ\����ٗ�����Ȕ�}ռ�,���Ÿ:�ǯ��V: K/��?1�yK5�Lxh�3Sxὂ�$�i*��{{�F�.o�֘zO�+�u�ye����\`�%�~�8�Z_F�ʨ��9i��g�U��Z�:Ѐ�6�(�PS����D��:�Χ�V1X�)"Y�k�a���r�[	���&,,�O�ṫ^�U�R�@n��}'jY���[�x�0��'x��Hn�<@ɪ��d�n+&�D�g�<Ζ��r� �(��˴x���;HkU��w��K�� �Yo��H
�n"�0T�O`G߳�*�i��
Ж�Nj�;�_�^���i_!�x��2���(\ n�ޏ��Ѫi�ȸL�8���3�����Wr+b�B�_�՚)ٖ�&��n<|�0B�`ˉ)X�D� I"�}��X�mvn�>�
6��F?��35q�M8G�=�̗��Dw}�LL%��R�5Q�R��}�آ�����5C��������F׼���̪D�Z��U���\XN����{��:� f)�WY�2���Y��o�˼6�wv"u�Zj2�;��=��L�xg�k_�r_ ����k8�/�8�V��&�f^���ب߿5�#O(k�_L8������n�wї�v��+~1II:��k���>;l��X�|��/7,�&-�	���j�R>�uf.[-����n1j�I�#��<�v4�;ձ�jN^L+` ��EG�!-�X�a��ϝ�m���aLrUl�?ፕ�G�Tp�].��w�x�	q�~��MH�����u��R�9h�����wDn"�=6d)�W�%��G�*�({��a+v9��'qWρ
]���!���ꮲa�HZ�:t+�o���9�"�M��WN�F�sgL8�Z?����ɩ�� 
��.{�Y"
�wv�Y}���b��A)ĉ~��џ�.��q3XpnY�z6��ʴm����g��\𖑿i4��Q����2md���R+��ao�%bE�.	���2�c�%EWI�\��K�Z����n��fdlh[I#%�����,�ÎB<y71Ur���Θ-{�ue�i&AI�W�m��8����Ҷ2+PA�Rx��v89�S\E���+Z�I�u{��N�C���l�Z�>�:;P��u�a�Ɵi�rΚ�F�9 �:����}R���z�nȢ�sT�D4��IA�i� ���4�$2�y"F�A���}�����~2�?�2](��ZHfڗ0���>�����l����*\A79�1=���`Pd�V�;a�[Qp&7��^��X�¦]���q]W��z�IR���s��1eBfH$gϗ7��N��Yh�K��6gk3�OX5�r�}�j~p~�$�f�LԾ���6˵��\��Tw<l����3{s֌�9xxe�
Щ���ί��}�"UN{���}�`Dk͠?��P�;�T}@�u"�vf/X��>ma�~`��N Y/���Bz�Lg�M-���ڻ;HU{ѳ��
h�Js��n��Lm�v�uLD�^�����X�c�y]��xfl�S�fF{5���^Qg���$t���߇%�*x�F� <�t��9OwD�C��{�8�k��yzN]Xi��2r[�Wͻ��?6ג������zV-�Fm��s�;��t��	�^ݼ�;���k�Y�o��: '��ɝ�}����4J�{���~cq\�Y�w`m�[cI�|j��X��=O�).Me�����=�,jǀ������Y�=E�� }{�1J,��2�U�}�ei���i3��?>����e��r9皇i̅r��)��a��Y2L�&+ׇ˵L����$Up��)&/�lYN���{�ʐ!&'�8Ta��..����i������w��!�.��P�?��\�<hǌ��GCS ���d����Uo[�k>/�[8D�#NM�����f�V�g�S�*b0+dg��&N��z�6b�S*�k�\�M������C۲���2ih{]����f�~�$А��
3��,�(Jx��Y��� '�?�d��\2&�;�Ai����Y�}��W�gJyF4�|j�
�<[�%R� -�v�<�X�B��X�nuյ��[� ��퐋?@H(�5΄�Y�]��uN��!��w8�n��`�{�=vb��!�=еK�Vi���)o��x�/��JY�͋��fnl��F���z���Tۨ�\�K�˽��v]hJ�8T���D�Fxx]���Y������i��M��0YA��>r���Xw#�I�a	�.~�����͝/�,�d���kV���ҝfk�k�����(�����?}���vEg+�kO�*��1�*}XŽs/[\�
I,����7��U ��-�v�?���W�mU-w�R��,����ȴ�D��z�z��;'�TA�S`�T�uJ*Z �5��Z�^�����aPE����ߡ~ئ�|Ru۹x�3:��>qK����p�e�Dro�S��-�
���X��\A�#�mz���g1�ᩋ��i�����qHsY�:����'E�Z!���Wq!����\}G�c�6�"B���6��ź0%�����CIz�3([.�0�t�{*?�"#c�N�W�����چm �@���X�M�f����萻���vՠ`�\fk�T=������DN�&)�K��"���/J�p/�������VeM����������siK܎�%�q�Z�\U�q��4uxN�H�>X�E��9�{�"^��U��=�v�1��2��,<�������YR.T���D��%m��wP��]1[��z}Z��F�ځ}̘+�DΖ[q�q��&�7�.r��n_�^c���ā>������ZO��bNm/`��ʐ���+־�ch�� ���V+�����\<%�u5u��E��E
�w%�U�j
�S�$t1�I���$�n��D��y�}��i�8���Cv�N�X�^�vN�s"�+9G�B��̔��Hm7��'�o'ˎ����[��;)��l�P>���>�O����QA��|9C7��]k��al�f?�$���WjM'�}.������U�˟�.VQ�Q�p�K�h�f�����{�5��a��`U� �^�05A	���3t峳:g�V�	Q�k:X8pz �}���2K�]jf��+_����;%���=|� M�L��Q=)��ŝ�����x��.wL�t棕X�Y�&5�Q?�ʿ®3����h)`�u�Dba�)�|�:mvs3�G�z�qV�[���Z�*=���M�b�1�;P/v����'�YDQ.�9�Xk�i.��?z�w�G���KR%��C߸#\	�"�M�K�]:��ln8�7'[x{mn����hubj�&��Azy�@ɋV�5�<��MZ�C�i����&�I�W����V�/�V-��������:	��"[����jn`�1
PG�N�P?�?��ھ�9���N�lJ�s�"H~TV��؈�)��vs20���2ݳ���r�B��BC�WѢ�wj���	v�EEJ�6a�M�L�����|`%�l[K�zP�vP�9Y�#!A5���&�6uT�<��R�-X�K�
_��y{���x�E%N�?I���?s�o0	��|��,��/����m�[��ӊ�R��k;��n�B�Co�����$ϙL��\+�N�c�N����R{η�p���r9�(��P߾�J��CY,bd������WXK�eo<���sG�(<G���ϑOf���.XF�~�VYZ�nm]Hf�A{��,��O�c}�G��B^o��1����T�\
�8�V���#r/�l	��Њ��߫X����Wv���>�
�~.ӫ�	~@Lb�7�H�B���I�}���3D�B��Ν.Z
��:	}h�XW=T���!v�u���b�K.NC'��8���A���Lհ�¬Ra���:["����j<�S�cM��5dzp���K��;{bB��l��7h�u?����V䱆�)xnK�u��mF���;��W�LX���$:0e���K�N.b|.UL���J�AJ��N���d��;�XA���5����vz�/|�@�]C��c0tHIw����Ο0P�^����.����PZ@��:�zYv��6|�u:6g��(�Aq�ʨ��	ad�r$S+/ـ��ڪW}�VЎ
�����]h�4��h���)��w*虨+��v�:��i�O]�OH[~��7����cQg�DSsi�a����Q��k�-��5�ڦ�TidӃ��߹������LD���ߑ+97,F��	�L ~R�M����\L��=U�yEem8���qg*GS��B�E��!��+�����WC��d�Y�~�^�E4�;������f5��'$�Zܥ�'�Ҹi��ė�_ө��9�_"&��f���:��_*(��P������AnZm���xw�R��t�$�2���?��5擥Cg�P)�Q��<'BW-�F%�g�q��6RR�
`��y$������.X�EY�I�<��`����Ѓ=B<����cD=W_k��IzP�o�.Tԇ5��Sе/���s$�CÇ��P���I�����`y����5���=�G�� :k\!$ِ�� d�2�f��E�V�\�۸QP�Z�O�r[t.�pMiK�6��Q,4&��)9�]�Ȝ�*�m�@�����O�ȼ�!j#��G	f8��)j�;1��l��Gi��r�N�ҔA�Fv?3��	�"EJ�{���$C
+a�q�����?�iķ���&T��]OH��mҝ��^�ǭ$������c��ڧT��	6XY�ZG[y�J�bu�4�/���S�
��E�k�/Q������o��I���孈>�UAӁ�W�O�:W<<1��ơ��^�{�-W�Szi��
Xl���/��W�"A���*<:)6�?PF�D�8R[-ȵ·z��J��t}�c��n�ʆ���䭀�`2��d|�T��	f\H�۱I
�-{LSL�K�q ��ϒp��6�������:�&P� ��AS�}eV���e������1t�]��CD$��S~� a\��B{��v8=D1��a#!*K���k���JH�?�2-�0�hƇ�iEP�4$꣰���bA��5�tX?�k'׊3�!�GVi�{\6q3/Έ��=�w4�%������!$k���_4�g�m�2����XF�r(�)ߧ����/�АS�:V9��������M.��ϒ�����ܥ?T�������+�V/������E���8mdI� �ln�f��VC(Q�ÛU=_�(�i����Lu�+.َ8��_�ڞT�qߩ�r���C�e�Z�̘�S�1~B#��_Iy�!���{�Wg�"�")��c�������]��1������j	���h\l�)n�a�)��'�by���*93!�ys�Q�b��(Fh9\+8cxT�ώnR8���{���h%���w�q7�_Ub�h���L	4 ��=��?�F�c��x]���7R�{��t2'���W���9�El?�+d���B�����S��˶-ǮP�J8�q*���HN�M6��yɮ$Q�6X�Z,Wĕ^�O]d��24��o�L��l�������֏	!�z�a��t�iS����㝾U'U��t+O���y�'��oH�J^=@o�0�kf����I��҈F�H�d�k��E��T^���h��	���9"�׵q�(ԩH6�;lmkP���Yu@�]c�J@�� tV�Q|��rx�=�w3�c��^�i�R$�y�O���bؤ�F��6owʦ�*����Ǳ��ͯM�X0b���J��_��*<����8n�=<?��+�n:��귐r����J�q�"�F'��"_��ݲ\;"�v��T�PWt>>*�Y"�ߍ����qE4��X+��l�����Q���ޓ�Ɖ
j�L-���l*+�iv�_U���8�}t���a�	[=�'( \�H�¥U��i�C�(h�A&, �e�$�p��U�nc�_mX��H� �����}�4f��	�a�Wt�	�f�@';��64�歊���l�劰��G��-R��b���D�'dq, y�ʾ�fK����RkR��~���6�/�qv^F��;����퇎Ȯ��@|�Є8�yY��ιT����\�r���U�SNC��zW6���eF����5��U$�I>A�WD�&~ �Ʒ7�,D�#��q+9�����NR�	������%�*,�I+�r)J^~�έ�]�I����h�D�	@[2���Co�Oq�T��/Ww1!9]�#E}ae�q��<�Z�J�?��-ɚ�$��oJ�\W��?�@%Г�8T&�/w���)rHJ�;�	�gB�ci�dB*�Z��y�qp{;r�0h�/��������������<4�y���aj����*���Gz�G?~5fA���d+�!\(:1�f��D3�J��(�o	�mA!֞H>�$w�O��/���M�_P�6��TXM�u�g��!o̽����&̆��c��#�'{�FC���dE;�g�e�����&����ݙ�Ƭ��/��K�~� d�X��9�S^VХĪ�ng>��1������{�;H��	�[PJ6��ꎆ��}��N��$���0�E�T`M�Ph��pG�Kp��3����%C��a�?�}^�-�$�U?��W-��n��Q=[Y�ެ��������0,�G�9�D���&��b�[���U��t��t>I"cC�S���0D
����K�t9�����D�>|�hH��	��	�f��1�-rq���y�A$E?M�K..z�Iǿ�}�
�M|�;��i��VG��4k=Px1�G��=��򒧒����xlۭ�f��S-d�#X�������Q��~##��q(�?.�ڴ��'R*|�lnP���s�d�S�����"W`�P)9�$����G��c��eN�/.r ��'���o0����b��!V�,C�̚���0��I|��SV���W��$�M�P��V橾���i/�ӶX>Ex�J7r5�����k�䊓Gn��(Or���������� .�ڰ��n�P#�.V[|ݻ�R�Y+��o�7m���Ί�{�c|d~�X��*Ti�mN�J�֎{�!�D[���������;��T�ش�	,d����g���\�B3]?�,�g2�~�C�p��qv���7�<���QҏyM'0�P��wV8W�yZd���y���9}�[��c��ܠ���Jy���tq��][��r] �>�8%���TVd��$e�N�@�}�&%S�Y�V��:2 7=7ۗ �A��&��T���4����H��/it��������b�R눜�u�B%��*�`	�LSo�T�Q:�uP�Ɍ��c�m9é��WMR�+�|)�NE�]_'L���0ik�l�XzR��$h�m
�����������Bܿ���m�5whM���*��;�~�[�YXY�]
[%�iqP��1�Y�_�&�U�x���h0K�'�_�<S��?��|�ulRy�ꡲ�!|��4� w�,{l�87��ٗ��w���JC��Vh�?�ۖ϶�~S;���$�Oը��>Q��U�2�<�����S��B]R]���O�d�P&^�n��1��G|g�rbm����'"a�gOn��0�a��R~���Ƨ��c��L����p���;��_ҷr���e+�p�|���hΘ� ��Q���6H���H�#��uĒ��v!};�?�3�1�I7�m���
���:Ћ�^�hf�W\r�x�8��8�n}�b�����(�c�pq��gw�����;8���Y�_ ���R���:ɩX��扂�ڑѐ��/�����9����U8R6Յ ?S|��-x��S ���o1V�r�e��Er��C�7qc2r@a������4h�w��n����d�"�Î�a,����������д:D޾,��	YM�{#0���!�Kt������b^��	���<ù�J,9�&{O&�	P]{��MEn�8?���`.��[i+�*���%��K�\H�Sv��b�z��4�	r�1-%&t ���ه!`�^N�TҸ�%�s׮;P�/��.�2��r.l���E=PY�mv�HT|	zcW��f��^��9Y��/0S��Ka�	�m�g_i>̰���I���d�v!�#��L���זeD]'撝gs�ΆN]m���kjg�ޤ�{`_�gs��������'���q큁V]�S��R�'4��(g���Fk���8}����1��d��5ɶ�d�C}�s�����=�J�� ������ˮ(4���Ќ����{�0�Ts.�&#�̆��ո�7ҹ�����e�zJd�!:�%��IZe 邅Ř|����J ��� ��[�M�j�Z��?g`�[�����_:H�-�w�	��M�ದ7�t_�vW)�����|L�#���m�M��c 	�ܴ���j��{~)U�',e��3'ŋ楩��긫��j�F���W�|�S'hz8����EU2@�?I渝K��k\<�̴m�H�P���{��H �ᗍ�fĉ+��(�ol��N�ȗ��"l�I'���N^È��OkquվR��O.4�q藳˻&sETr��B�s����8f�|���'*t�9���P�քϊy(�4�' pe�܎+��"E*��^���(K�
��~����D3�>�vt=��Wi>�Tzy����@8��q��lO{�Y�ݩ�Y�}&O^�(W
ɪ0�t[�Rb���+5�$	`��Nh{��QůP ���}�HfW|����HX"�/�]Z���/KE21LT9̗w�SG +�����9ѧ�tfχ�_�g?*��!��kЎ�ݞr�^Y7�p?��O-��7h�r�xl��EWq#���0��/�߲��/B"�_��p�e$�v�:d$x�[�� V��6�&��5��rD���@��Z�]S�
�-u��I�AIv�J�*Z�G�wő2b���5�q�U��s���O�9��<���)�\Â��*v��d	�g��#�׃�\{0�_I4��q��ӒD�z.�!�l��YF&6�LA�#@�H�Fx�~�@��eU84��<z�h�%� ���=f,^r$�A���'�d������5o S~��3�`�*q�c�r���\�ґ�g	2A@��F]��9ua�!��eL�A�P�bi�!�<#m,������9j]�l������w:럱�E,$�<��K��+�8���V����:*���/�e�[i��V�v]�`L�v-� ��y�	.v��B��ip5J`�9��K�|����I�D �����[{�p!��(�/Ф*d��\DG�� ��1M�pF��x��u�w�O	�5�-�<h6�X!cvckW.�ͤ��Mɒ)�;��3]n{�?^�:�j3���p��4�
g �6,���O�_�.~�ސx<6kF6V�:u�Z҇+�#1�q�}��a]��!��O�"N���]A�R��b��oet�������7q/�,��c����_1�I�
�fK(��Q\:��<nHc�Sj%�ԑK������;��?���3N�H#���|�<|&I��UY����B)~���+ԯ�1I�T֠��Ka��IO�]��^x}��߫�/ ������-�2i��
蹁Ϧ�B4-{�JٻҡYu��&=�ôE���֛���ï�5�[@F�L���y;�[ah��<�|h���A������f���|��Ѓ�`Y���y���h��"����6�MdS�p��,��!:�Y��B���e��O�I�Wf��T	ۑ�u�����9�L���@�ە��Ot�E�e��g������x�Hѩ��Hk>�p��>��u��?�mp��w�7%0�(S�fU5��9��֎o��ʁ̫��r%���Ԫw�����K�v���JnIt$dsI�zÝ�O|�Š-u�������R�A;���T���YH�����M��2x�?�:���*�Ȧ�[������>��s����z���l��!Z��O};��ul�5U�!}�A��,���Bg<���8�1�Y�zr�/o�n��u�E�Yk�ܵ
n�ڛ,i{����(�X�Ss$`_@�~�!b+�9n�0�������D+���q���V���%���}<<�"!��eh֣Ua��P�R�>5%�SJB���S���s���*ꭲ�/ъ��c��=�/(P�R�B���]ToB�VPt,'��|>��~��ma��
ŧ�J�)��e��CR�9�JO���Ztf��L�7�2?eO��|��T.7�
��iN���F����Q���`'�
�@=���˥.`�
�NgJ�*�M�s��+���š����Ҁ�f:�8+�,;k겏��2�����1T4�P
̂�:�!�b��{F,`��F1$��Z��,�##B#�uk��j)�y��i{���p6��,�(J�