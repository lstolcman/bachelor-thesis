��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J�-�4ϼA�IŠ��#�U�(�f���+�p-Hv"�-L��wUoV�5�󷹿1��4��[c��i�>�cű�A��&;"��+p���N�'�p��gMG��6l�7ֲ@eo2;��5��_<\zڪ:C�EwZ��6�&x��Lq?��n]�9⪎�o�PE�G�k�ڑ�O��f�;�̍Y"�)ߞ�m̷����#.��؜)�	NY=j��R��#o(��2W{���,Z	�H��Qkٝ1���0p��z����9!�Zls��#X__d���(�_��I�^���-K1rS}ݐ�UGr�ܲ�F��6�c�W������!�U���H�4�A�`�QJ����gy��&��^lqʵ(�ڎ>I��6qTr��0@�j���#A�u\k�����$o��v�V�-
����y�_)� \��0�.��4�;q�z��7w��qs�>���R�q�-}�ei�����$����t����$��F�V`�������A@��nR7�������ɫV���3	$fld�u��-��c��*��PZ�6[^&�$>1���SIF�� 
t����G
ޡ�yS�Z�X�M�.=�?��Z��@�N-?9�k��ЊVP�:�]-���.�����^��&o���Ǧ�f�Ubh�����s��u����94��0;M�G���(�-�J��}I��*޺\� XO)�:��5�r����D���Ōv�[E|%P:?��=A��#/3Mi?"�o��G��f_Q:��Zw)��d,1�a��ގ^�V�D�A�f����c��W'�D�������=�t����(]O����a!�w"#a}���Ǭ ����0��Q��/:�!��&'͑��"�V��|��.!Rk��s�K��FF1z��3�/}.j�W�o׊f.��aS�h��� 7H�{����g��U�����KP�d�>�F����:!��U�+H1�2��ON���.���j ��TX����7������zẐ2���md���l�C�Lb@���=T�_˦�buf� �$ѥ�� =�"͗Y�m�6_��P�h����JZB��]�NAbচ��֨�T0X����i�^K�̐$���]F8+Q�?9�
Mig���G(��ٖ�X�+�N�q��S�#����>_1"�=���Qh��w��ì�;~�4���I���|�/0�6$��@XS�a���/����3�v����׎���N$��bF9tl�ӜZ�k�`���|�芪�����]¢V�.!I`U`�o���a�Z��NMȢ_���m�-����髩"<�x(�AR�:<	��(��u;��6?�\���&t߄��{x���Wj�t�jcP�G��P>��_�/,�{�c3F���Ys3�1�1��u�,��o�h:WI�]�Wz���|>�z���,�;y6��V�ݓa��v"�{��3Mc^f2c�Ɏ���`�t
�W�c �P ^ �٠���pH%G�3P/0��k�5R�3a�q&{���r�=���?X��=vB!:U�j��j��u�	�����C����^^\��VA�LE����XS�,�j8��"�GE��b�X����@\=�ؖd��IZb��N�6�W}N�:����\K!��Ƣ��%4��0�r�Zl7�����^�߽$!w�°�42��[r���g�AV�l���8
Rp���Lu�5��|�ǿ�μ�3�:��`8��7zW=�Վ�q�"{�{H��m��yd��'PGY@�Qr��ʀ��a��Z�,d��g�����-0� ���eN<�H�[�9�P��T}��_Z$N$� 0�����*�����5Wm���#�'��mA�썁o7��3���8��r�6=�_U'Ǜ.�#�����gP�r=0���lM8�=/1�N���M�)�z	̣�衮�n;
�nX�XՎ��kwjG�RI�~��Ԯ�t����S~����8�<���9�'�VA�I�G�2��<{�Z���OA���93���u��κ�xl���Sd�<�nA�!#���6�"V������1!؟���b���)��0.#P$	,��HsZ��I�ŦW�2����qI'�9�����kc�)̇p��MQ@{`�dY :b�E�.۷��P#��En:jQ��[��� xbR���X.Na��䭾�ѫ��GIG�7��V[^���v��w�Jg�o��GB{%%x�mB}�P�ߊ��h��w"�U���s}ꬷA�6\Ī��kſ�p���I��X���,� q����>pO	2�>E��]&Zv
��AkE�� �1T�V�*3R3�fpߑ�D�F�ݜ�F������琮;��g���"�vi����E��Ȕ�~WrE�R�C�TTo;�V�%� � ��܂O"G~u��4�1Baˍ]%�\x4�9��S	��H6�+�Z>Ϣ�B��V�yb�� �n�Z�u�9i�)�'�������bk��H��G��$#6�w cl{Yθҩr��p�o*O��b
#�2D��BU��ܜ����C(lݎ5��kbk��J��'J5�h����d��TI�VD��&��� /���|��Hp�@௏���7�����.�>���Ok����;2�C���j��e
�k�p�P�P0�#	���`�:����V����9�j(m�N�/��c
j�h���R�k���k /��z���@@�^���P�R��2��Y�Uz�{�yڕ�M�Sp����Yӷ?���H�w�8�/�z���y7C�=�#'�k�<�F�����9r���/��e���ޯ�u�z"��E U�$W&��m����H����_��7�0
h�����{�'�1H�k������e��G��AɊQ7��a���-)�:���+Q��U�[2�I[�d30�Ww��S�\�Ӧ�Dh���1mP~�-����D�C����X˫�����tJ�΍q>=�x����/�⨥�C��A(�]��J]t�H��9��D�nʧV����Hm]-B���OJ4��І��]��5�u}���M�l>�u�N]���'�h}	�%�ʼ?yS��7����BP(���{�
W<�nև��ګ��w�G��o)���v]�5b�����L���b+x?�=KP��O<.�U�`�}}�$�$Z%��w��L��'x�POC��_4u0�YPt��l��k��08�g�Q~Em��H�	������'�r70�J�Q��!b�|�ɟ���i �pZz ��P3�Ϻ�����Ն�i��A˄��ƅ�[����������V�i ���)���R�8:{>P�gQ���g+2����V�H�bK'm�0�l<�U��h���u���1F�i�㨍SN�V`���X�?��<�q��#h�1��yBO�{�nPZ��wg^ӮR~�vB�xd �� �$Ű��a� �Fr�Wm�F$��c>_��^��7�af�vOҞ���H�Z�Qn?�t�z�{��m�pr+�SD+7�	�
a�n�4VEoXpJ�_=�9��r_�����~����N�j�(�b���~�H�>��Rw��s��>��S�rrq�<f`�R�����{>7�Q��=��C-: h�7!�HEbv�j?��l�Փ��;�g�y�#�&�~�+]۠\�/��1aw��@|��H+C�B�0��0L�⡙�< �?��UU����կ	fA��3O�+=v�D����?�Gz�RLNO�'���� F���S۹�h5��	�ϳ�8�S�kl�z�h5��n���rvPC��f	���l g /���dr�U�^�C(*�5�R��j`�0��&�=���6�����e'��1)����'���wi�77v�^ھ��k90i����Ƒ���LM,�"(���&�����F�oI^�\�"�8����;	�;��Ƞ,�B�~d��FJ�qyQcP�
�@�S��}��.l����w�$kAC�N��w�T,9� ��>��~�.��x�u�jf�L���I��P�]�|y��p�b��P���6�u#밷��Єk.��������4��;��/��A:�>O��'��ػ�zᝠkg���/�
'�]ȁ�g���;j���^۟2}��y%ka�s��AgG���Bf݆W���#�3���m
�<vTv�G�3-��k�i�O.�I$�uA㬬L�4� eA	+����5D���J������%i�s	��X(u�ȇ�ٲ񶒏���W�/�X(F�VmH?�s��R�Qށ?���WƟ�C䧤������Z�{� ҵ�{M��=!��9|@)����.�]�dm���'��ܷ�V���Sw,��ϓiB���?@+t�D5�>Ce�P72OK���[�������&��ܓ�bI�Lt'����>�P��� �Y$;���_��?1\l��Y�ך�<�vf֜�_A��^N���d[}��d�Y����h>6ʶ�d���`�1��TwN��F��g�A�y,D�]���p���=��eXI�����R�G�4؁�-8�Lx�LqO�[��N�Ud:�A��Y�X#�Vʆ�k�� ���'�^�٘�:�kS�rF�1Ox�ca�(�O����29%�zy��,/�I���PH�j�����"������9g�7
yt�B�]���d�9�n��=����1��r�<�,t���r�9��o�YK7c��c�������������;��ՋY��
o���� ĚD}]��Ȑ{��7䟨T��%��S�S�G�^��7����0�IF!!�v��$_�@��ِF;��H��։�;���r��7U�����ZqV���2��x��EbDj�H�v��WL_!��8�SҩI�<�:c�O�G�� �|L��P�V�kOsʚ��=�^0����%׳/rt9�@u�N�vd��q����l�
U�F���cS�2L2;3�`�� ��[+�͓�Iw����`����[9uдNlɚ��¸K�}��E�mCdH�txqW4\�/i��Z9���n5 �)W(����u���m, �St�����}&�(!�߲��!�-)PP�/H ^^�7n��*���p����� �r q|��?U� �ǳ���K�9/g�fܝ��5������ZN3�E�ϥDɴ�)J�p�
�מ散rr��Mf���<E;fK��0����m���x�h�lGi>	%qe�Z�ߵ�s�� g�FI:W���8)�d��q2�X���b^��O�<�T�]�m�]t\���Pn�GU4c��*W�	�,�?[�.�J�u/�yW"ŉoھ6��\�Ѣh78U�s��nU���F�7��J�A���#S'*7�?�B@_�_����7��lP�6����@K��8���ְW�1�,}J��_��R�ٿK���k��׊Z+~��d��Ť�袇���=]�^z���Ӝd��i�����?w���3s��
+~��$v�s+���ƙ)k,֞�_!�ML.у����_V�gWꅰ�=�o�V)g�7E���*��'�\����Q�u����X������+u"��I�t���;4Y���gԛi>�4Rf%X�\�T3��3�
Ȅ��ՏV��1�/d�osB,��v�+nN�5��+m��(�"������r�T��3����g�